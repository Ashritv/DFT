module vorca (clk, i_reset_, i_sw_init, i_addr, i_wr_strb, 
 i_wr_data, i_rd_strb, o_rd_data, o_ack, o_err_ack, o_spare_config, 
 o_adj_config, o_dbg_config, i_revision_config, i_spare_config, 
 i_hb_sup, i_hisbuf0_0, i_hisbuf1_0, 
 i_hisbuf2_0, i_hisbuf3_0, 
 i_hisbuf0_1, i_hisbuf1_1, 
 i_hisbuf2_1, i_hisbuf3_1, 
 i_hisbuf0_2, i_hisbuf1_2, 
 i_hisbuf2_2, i_hisbuf3_2, 
 i_hisbuf0_3, i_hisbuf1_3, 
 i_hisbuf2_3, i_hisbuf3_3, 
 i_hisbuf0_4, i_hisbuf1_4, 
 i_hisbuf2_4, i_hisbuf3_4, 
 i_hisbuf0_5, i_hisbuf1_5, 
 i_hisbuf2_5, i_hisbuf3_5, 
 i_hisbuf0_6, i_hisbuf1_6, 
 i_hisbuf2_6, i_hisbuf3_6, 
 i_hisbuf0_7, i_hisbuf1_7, 
 i_hisbuf2_7, i_hisbuf3_7, i_agg_su_count_a, 
 o_reg_written, o_reg_read, o_reg_wr_data, o_reg_addr, scan_iso_or, 
 test_se, scan_iso_or1, scan_iso_or2, scan_iso_or3, scan_iso_or4, 
 scan_iso_or5, scan_iso_or6, scan_iso_or7, scan_iso_or8, scan_iso_or9, 
 test_si1, test_so1, scan_enable, raw_scan_en );
  input [7:0] i_addr;
  input [31:0] i_wr_data;
  output [31:0] o_rd_data;
  output [31:0] o_spare_config;
  output [15:0] o_adj_config;
  output [0:0] o_dbg_config;
  input [7:0] i_revision_config;
  input [31:0] i_spare_config;
  input [2:0] i_hb_sup;
  input [23:0] i_hisbuf0_0;
  input [23:0] i_hisbuf1_0;
  input [31:0] i_hisbuf2_0;
  input [27:0] i_hisbuf3_0;
  input [23:0] i_hisbuf0_1;
  input [23:0] i_hisbuf1_1;
  input [31:0] i_hisbuf2_1;
  input [27:0] i_hisbuf3_1;
  input [23:0] i_hisbuf0_2;
  input [23:0] i_hisbuf1_2;
  input [31:0] i_hisbuf2_2;
  input [27:0] i_hisbuf3_2;
  input [23:0] i_hisbuf0_3;
  input [23:0] i_hisbuf1_3;
  input [31:0] i_hisbuf2_3;
  input [27:0] i_hisbuf3_3;
  input [23:0] i_hisbuf0_4;
  input [23:0] i_hisbuf1_4;
  input [31:0] i_hisbuf2_4;
  input [27:0] i_hisbuf3_4;
  input [23:0] i_hisbuf0_5;
  input [23:0] i_hisbuf1_5;
  input [31:0] i_hisbuf2_5;
  input [27:0] i_hisbuf3_5;
  input [23:0] i_hisbuf0_6;
  input [23:0] i_hisbuf1_6;
  input [31:0] i_hisbuf2_6;
  input [27:0] i_hisbuf3_6;
  input [23:0] i_hisbuf0_7;
  input [23:0] i_hisbuf1_7;
  input [31:0] i_hisbuf2_7;
  input [27:0] i_hisbuf3_7;
  input [31:0] i_agg_su_count_a;
  output [31:0] o_reg_wr_data;
  output [7:0] o_reg_addr;
  input clk, i_reset_, i_sw_init, i_wr_strb, i_rd_strb, test_se, test_si1,
 scan_enable, raw_scan_en;
  output o_ack, o_err_ack, o_reg_written, o_reg_read, scan_iso_or,
 scan_iso_or1, scan_iso_or2, scan_iso_or3, scan_iso_or4, scan_iso_or5,
 scan_iso_or6, scan_iso_or7, scan_iso_or8, scan_iso_or9, test_so1;
  wire N468, n468, n265, N469, n469, n266, n267, n268, n269, n670, n671,
 n672, n673, N470, n470, n674, f_err_ack, N471, n471, n675, N472, n472,
 n676, N473, n473, n270, n677, N474, n474, n271, n678, N475, n475,
 n272, n679, N476, n476, n273, N477, n477, n274, N478, n478, n275,
 N479, n479, n276, n277, n278, n279, n680, n681, n682, n683, N480,
 n480, n684, N481, n481, n685, N482, n482, n686, N483, n483, n280,
 n687, N484, n484, n281, n688, N485, n485, n282, n689, n486, n283,
 n487, n284, n488, n285, n489, n286, n287, n288, n289, n690, n691,
 n692, n693, n490, n694, n491, n695, n492, n696, n493, n290, n697,
 n494, n291, n698, n495, n292, n699, n496, n293, n497, n294, n498,
 n295, n499, n296, n297, n298, n299, net121977, net121972, n700, n701,
 n702, n703, n500, n704, n501, n705, n502, n706, n503, n300, n707,
 n504, n301, n708, n505, n302, n709, n506, n303, n507, n304, n508,
 n305, n509, n306, n307, n308, n309, n710, n711, n712, n713, n510,
 n714, n511, n715, n512, n716, n513, n310, n717, n514, n311, n718,
 n515, n312, n719, n516, n313, n517, n314, n518, n315, n519, n316,
 n317, n318, n319, n720, n721, n722, n723, n520, n724, n521, n725,
 n522, n726, n523, n320, n727, n524, n321, n728, n525, n322, n729,
 n526, n323, n527, n324, n528, n325, n529, n326, n327, n328, n329,
 n126, n730, n127, n128, n732, n129, n733, n530, n734, n531, n735,
 n532, n736, n533, n330, n737, n534, n331, n738, n535, n332, n739,
 n536, n333, n130, n537, n334, n131, n538, n335, n132, n539, n336,
 n133, n337, n134, n338, n135, n339, n136, n740, n137, n741, n138,
 n742, n139, n743, n540, n744, n541, n745, n542, n746, n543, n340,
 n747, n544, n341, n748, n545, n749, n546, n343, n140, n547, n344,
 n141, n548, n345, n142, n549, n346, n143, n347, n144, n348, n145,
 n349, n146, n750, n147, n751, n148, n752, n149, n753, n550, n754,
 n551, n755, n552, n756, n553, n350, net121966, n757, n554, n351, n758,
 n555, n352, n759, n556, n353, n150, n557, n354, n151, n558, n355,
 n152, n559, n356, n153, n357, n154, n358, n155, n359, n156, n760,
 n157, n761, n158, n762, n159, n763, n560, n764, n561, n765, n562,
 n766, n563, n360, n767, n564, n361, n768, n565, n362, n769, n566,
 n363, n160, n567, n364, n161, n568, n365, n162, n569, n366, n163,
 n367, n164, n368, n165, n369, n166, n770, n167, n771, n168, n772,
 n169, n773, n570, n774, n571, n775, n572, n776, n573, n370, n777,
 n574, n371, n778, n575, n372, n779, n576, n373, n170, n577, n374,
 n171, n578, n375, n172, n579, n376, n173, n377, n174, n378, n175,
 n379, n176, n780, n177, n781, n178, n782, n179, n783, n580, n784,
 n581, n785, n582, n786, n583, n380, n787, n584, n381, n788, n585,
 n382, n789, n586, n383, n180, n587, n384, n181, n588, n385, n182,
 n589, n386, n183, n387, n184, n388, n185, n389, n186, n790, n187,
 n791, n188, n792, n189, n793, n590, n794, n591, n795, n592, n796,
 n593, n390, n797, n594, n391, w_load_spare_config, n798, n595, n392,
 n799, n596, n393, n190, n597, n394, n191, n598, n395, n192, n599,
 n396, n193, n397, n194, n398, n195, n399, n196, n197, n198, n199,
 w_load_dbg_config, n800, n801, n802, n803, n600, n804, n601, n805,
 n602, n806, n603, n400, n807, n604, n401, n808, n605, n402, n809,
 n200, n606, n403, n201, n607, n404, n202, n608, N405, n405, n203,
 n609, N406, n406, n204, N407, n407, n205, N408, n408, n206, N409,
 n409, n810, n207, n811, n208, n812, n209, n813, n610, n814, n611,
 n815, n612, n816, n613, N410, n410, n817, n614, n411, n818, n615,
 n412, n819, n616, n413, n210, n617, n414, n211, n618, n415, n212,
 n619, n416, n213, n417, n214, n418, n215, n419, n216, n820, n217,
 n821, n218, n822, n219, n823, n620, n824, n621, n825, n622, n826,
 n623, N420, n420, n827, n624, N421, n421, n828, n625, N422, n422,
 n829, n626, N423, n423, n220, w_load_adj_config, n627, N424, n424,
 n221, n628, N425, n425, n222, n629, N426, n426, n223, N427, n427,
 n224, N428, n428, n225, N429, n429, n226, n830, n227, n831, n228,
 n832, n229, n833, n630, n834, n631, n835, n632, n836, n_write, n633,
 N430, n430, n837, n634, N431, n431, n838, n635, N432, n432, n839,
 n636, N433, n433, n230, n637, N434, n434, n231, n638, N435, n435,
 n232, n639, N436, n436, n233, N437, n437, n234, N438, n438, n235,
 N439, n439, n236, n840, n237, n841, n238, n842, n239, n843, n640,
 f_ack, n844, n641, n845, n642, n846, n643, N440, n440, n847, n644,
 N441, n441, n848, n645, N442, n442, n849, n646, N443, n443, n240,
 n647, N444, n444, n241, n648, N445, n445, n242, n649, N446, n446,
 n243, N447, n447, n244, N448, n448, n245, N449, n449, n246, n850,
 n247, n851, n248, n852, n249, n853, n650, n854, n651, n855, n652,
 n856, n653, N450, n450, n857, n654, N451, n451, n655, N452, n452,
 n859, n656, N453, n453, n250, n657, N454, n454, n251, n658, N455,
 n455, n252, n659, N456, n456, n253, N457, n457, n254, N458, n458,
 n255, N459, n459, n256, n860, n257, n861, n258, n862, n259, n863,
 n660, n661, n662, n663, N460, n460, n664, N461, n461, n665, N462,
 n462, n666, N463, n463, n260, n667, N464, n464, n261, n668, N465,
 n465, n262, n669, N466, n466, n263, N467, n467, n264,
 o_reg_addr_reg_1__scan_iso_or_n, o_reg_addr_reg_0__scan_iso_or_n,
 n_94_, n_95_, n_96_, n_97_, n_98_, n_99_, n_100_, n_101_, n_102_,
 n_103_, n_104_, n_105_, n_106_, n_107_, n_108_, n_109_, n_110_,
 n_111_, n_112_, n_113_, n_114_, n_116_, n_117_, n_118_, n_119_,
 n132_inv, n395_inv, n500_inv, n353_inv, n188_inv, n199_inv, n343_inv,  
 n363_inv, n777_inv, n787_inv, n797_inv, n808_inv, n822_inv, n856_inv,
 n_120_, n_121_, n_122_, n_123_, n_124_, n_125_, n1;
  wire [31:0] f32_mux_0_data;
  wire [31:0] f32_mux_1_data;
  wire [2:0] f_state;

  SDFFRX1 f_state_reg_0_ ( .D(N405), .SI(f_err_ack), .SE(scan_enable), .CK(clk), .RN(n860), .Q(f_state[0]) );
  SDFFRX1 f_state_reg_1_ ( .D(N406), .SI(f_state[0]), .SE(scan_enable), .CK(clk), .RN(n128), .Q(f_state[1]) );
  SDFFRX1 f_state_reg_2_ ( .D(N407), .SI(f_state[1]), .SE(scan_enable), .CK(clk), .RN(n129), .Q(f_state[2]) );
  SDFFRX1 f_ack_reg ( .D(N408), .SI(f32_mux_1_data[31]), .SE(scan_enable), .CK(clk), .RN(n128), .Q(f_ack) );
  SDFFRX1 n_write_reg ( .D(n842), .SI(f_state[2]), .SE(scan_enable), .CK(clk), .RN(n129), .Q(n_write) );
  SDFFRX1 o_reg_addr_reg_7_ ( .D(i_addr[7]), .SI(o_reg_addr[6]), .SE(scan_enable), .CK(net121972), .RN(n128), .Q(o_reg_addr[7]) );
  SDFFRX1 o_reg_addr_reg_6_ ( .D(i_addr[6]), .SI(o_reg_addr[5]), .SE(scan_enable), .CK(net121972), .RN(n129), .Q(o_reg_addr[6]) );
  SDFFRX1 o_reg_addr_reg_5_ ( .D(i_addr[5]), .SI(o_reg_addr[4]), .SE(scan_enable), .CK(net121972), .RN(n128), .Q(o_reg_addr[5]) );
  SDFFRX1 o_reg_addr_reg_4_ ( .D(i_addr[4]), .SI(o_reg_addr[3]), .SE(scan_enable), .CK(net121972), .RN(n859), .Q(o_reg_addr[4]) );
  SDFFRX1 o_reg_addr_reg_3_ ( .D(i_addr[3]), .SI(o_reg_addr[2]), .SE(scan_enable), .CK(net121972), .RN(n859), .Q(o_reg_addr[3]) );
  SDFFRX1 o_reg_addr_reg_2_ ( .D(i_addr[2]), .SI(n862), .SE(scan_enable), .CK(net121972), .RN(n859), .Q(o_reg_addr[2]) );
  SDFFRX1 o_reg_addr_reg_1_ ( .D(i_addr[1]), .SI(n863), .SE(scan_enable), .CK(net121972), .RN(n859), .Q(n862) );
  SDFFRX1 o_reg_addr_reg_0_ ( .D(i_addr[0]), .SI(n_write), .SE(scan_enable), .CK(net121972), .RN(n859), .Q(n863) );
  SDFFRX1 f_err_ack_reg ( .D(N409), .SI(f_ack), .SE(scan_enable), .CK(clk), .RN(n859), .Q(f_err_ack) );
  SDFFRX1 f32_mux_1_data_reg_0_ ( .D(N454), .SI(f32_mux_0_data[31]), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_1_data[0]) );
  SDFFRX1 f32_mux_1_data_reg_1_ ( .D(N455), .SI(f32_mux_1_data[0]), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_1_data[1]) );
  SDFFRX1 f32_mux_1_data_reg_2_ ( .D(N456), .SI(f32_mux_1_data[1]), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_1_data[2]) );
  SDFFRX1 f32_mux_1_data_reg_3_ ( .D(N457), .SI(f32_mux_1_data[2]), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_1_data[3]) );
  SDFFRX1 f32_mux_1_data_reg_4_ ( .D(N458), .SI(f32_mux_1_data[3]), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_1_data[4]) );
  SDFFRX1 f32_mux_1_data_reg_5_ ( .D(N459), .SI(f32_mux_1_data[4]), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_1_data[5]) );
  SDFFRX1 f32_mux_1_data_reg_6_ ( .D(N460), .SI(f32_mux_1_data[5]), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_1_data[6]) );
  SDFFRX1 f32_mux_1_data_reg_7_ ( .D(N461), .SI(f32_mux_1_data[6]), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_1_data[7]) );
  SDFFRX1 f32_mux_1_data_reg_8_ ( .D(N462), .SI(f32_mux_1_data[7]), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_1_data[8]) );
  SDFFRX1 f32_mux_1_data_reg_9_ ( .D(N463), .SI(f32_mux_1_data[8]), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_1_data[9]) );
  SDFFRX1 f32_mux_1_data_reg_10_ ( .D(N464), .SI(f32_mux_1_data[9]), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_1_data[10]) );
  SDFFRX1 f32_mux_1_data_reg_11_ ( .D(N465), .SI(f32_mux_1_data[10]), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_1_data[11]) );
  SDFFRX1 f32_mux_1_data_reg_12_ ( .D(N466), .SI(f32_mux_1_data[11]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[12]) );
  SDFFRX1 f32_mux_1_data_reg_13_ ( .D(N467), .SI(f32_mux_1_data[12]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[13]) );
  SDFFRX1 f32_mux_1_data_reg_14_ ( .D(N468), .SI(f32_mux_1_data[13]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[14]) );
  SDFFRX1 f32_mux_1_data_reg_15_ ( .D(N469), .SI(f32_mux_1_data[14]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[15]) );
  SDFFRX1 f32_mux_1_data_reg_16_ ( .D(N470), .SI(f32_mux_1_data[15]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[16]) );
  SDFFRX1 f32_mux_1_data_reg_17_ ( .D(N471), .SI(f32_mux_1_data[16]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[17]) );
  SDFFRX1 f32_mux_1_data_reg_18_ ( .D(N472), .SI(f32_mux_1_data[17]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[18]) );
  SDFFRX1 f32_mux_1_data_reg_19_ ( .D(N473), .SI(f32_mux_1_data[18]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[19]) );
  SDFFRX1 f32_mux_1_data_reg_20_ ( .D(N474), .SI(f32_mux_1_data[19]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[20]) );
  SDFFRX1 f32_mux_1_data_reg_21_ ( .D(N475), .SI(f32_mux_1_data[20]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[21]) );
  SDFFRX1 f32_mux_1_data_reg_22_ ( .D(N476), .SI(f32_mux_1_data[21]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[22]) );
  SDFFRX1 f32_mux_1_data_reg_23_ ( .D(N477), .SI(f32_mux_1_data[22]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[23]) );
  SDFFRX1 f32_mux_1_data_reg_24_ ( .D(N478), .SI(f32_mux_1_data[23]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[24]) );
  SDFFRX1 f32_mux_1_data_reg_25_ ( .D(N479), .SI(f32_mux_1_data[24]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[25]) );
  SDFFRX1 f32_mux_1_data_reg_26_ ( .D(N480), .SI(f32_mux_1_data[25]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[26]) );
  SDFFRX1 f32_mux_1_data_reg_27_ ( .D(N481), .SI(f32_mux_1_data[26]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[27]) );
  SDFFRX1 f32_mux_1_data_reg_28_ ( .D(N482), .SI(f32_mux_1_data[27]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_1_data[28]) );
  SDFFRX1 f32_mux_1_data_reg_29_ ( .D(N483), .SI(f32_mux_1_data[28]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_1_data[29]) );
  SDFFRX1 f32_mux_1_data_reg_30_ ( .D(N484), .SI(f32_mux_1_data[29]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_1_data[30]) );
  SDFFRX1 f32_mux_1_data_reg_31_ ( .D(N485), .SI(f32_mux_1_data[30]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_1_data[31]) );
  SDFFRX1 o_reg_read_reg ( .D(N420), .SI(o_reg_addr[7]), .SE(scan_enable), .CK(clk), .RN(n861), .Q(o_reg_read) );
  SDFFRX1 f32_mux_0_data_reg_31_ ( .D(N453), .SI(f32_mux_0_data[30]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[31]) );
  SDFFRX1 f32_mux_0_data_reg_30_ ( .D(N452), .SI(f32_mux_0_data[29]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[30]) );
  SDFFRX1 f32_mux_0_data_reg_29_ ( .D(N451), .SI(f32_mux_0_data[28]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[29]) );
  SDFFRX1 f32_mux_0_data_reg_28_ ( .D(N450), .SI(f32_mux_0_data[27]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[28]) );
  SDFFRX1 f32_mux_0_data_reg_27_ ( .D(N449), .SI(f32_mux_0_data[26]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[27]) );
  SDFFRX1 f32_mux_0_data_reg_26_ ( .D(N448), .SI(f32_mux_0_data[25]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[26]) );
  SDFFRX1 f32_mux_0_data_reg_25_ ( .D(N447), .SI(f32_mux_0_data[24]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[25]) );
  SDFFRX1 f32_mux_0_data_reg_24_ ( .D(N446), .SI(f32_mux_0_data[23]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[24]) );
  SDFFRX1 f32_mux_0_data_reg_23_ ( .D(N445), .SI(f32_mux_0_data[22]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[23]) );
  SDFFRX1 f32_mux_0_data_reg_22_ ( .D(N444), .SI(f32_mux_0_data[21]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[22]) );
  SDFFRX1 f32_mux_0_data_reg_21_ ( .D(N443), .SI(f32_mux_0_data[20]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[21]) );
  SDFFRX1 f32_mux_0_data_reg_20_ ( .D(N442), .SI(f32_mux_0_data[19]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[20]) );
  SDFFRX1 f32_mux_0_data_reg_19_ ( .D(N441), .SI(f32_mux_0_data[18]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[19]) );
  SDFFRX1 f32_mux_0_data_reg_18_ ( .D(N440), .SI(f32_mux_0_data[17]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[18]) );
  SDFFRX1 f32_mux_0_data_reg_17_ ( .D(N439), .SI(f32_mux_0_data[16]), .SE(scan_enable), .CK(net121966), .RN(n128), .Q(f32_mux_0_data[17]) );
  SDFFRX1 f32_mux_0_data_reg_16_ ( .D(N438), .SI(f32_mux_0_data[15]), .SE(scan_enable), .CK(net121966), .RN(n129), .Q(f32_mux_0_data[16]) );
  SDFFRX1 f32_mux_0_data_reg_0_ ( .D(N422), .SI(n_94_), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_0_data[0]) );
  SDFFRX1 f32_mux_0_data_reg_1_ ( .D(N423), .SI(f32_mux_0_data[0]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_0_data[1]) );
  SDFFRX1 f32_mux_0_data_reg_2_ ( .D(N424), .SI(f32_mux_0_data[1]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[2]) );
  SDFFRX1 f32_mux_0_data_reg_3_ ( .D(N425), .SI(f32_mux_0_data[2]), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_0_data[3]) );
  SDFFRX1 f32_mux_0_data_reg_4_ ( .D(N426), .SI(f32_mux_0_data[3]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_0_data[4]) );
  SDFFRX1 f32_mux_0_data_reg_5_ ( .D(N427), .SI(f32_mux_0_data[4]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[5]) );
  SDFFRX1 f32_mux_0_data_reg_6_ ( .D(N428), .SI(f32_mux_0_data[5]), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_0_data[6]) );
  SDFFRX1 f32_mux_0_data_reg_7_ ( .D(N429), .SI(f32_mux_0_data[6]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_0_data[7]) );
  SDFFRX1 f32_mux_0_data_reg_8_ ( .D(N430), .SI(f32_mux_0_data[7]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[8]) );
  SDFFRX1 f32_mux_0_data_reg_9_ ( .D(N431), .SI(f32_mux_0_data[8]), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_0_data[9]) );
  SDFFRX1 f32_mux_0_data_reg_10_ ( .D(N432), .SI(f32_mux_0_data[9]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_0_data[10]) );
  SDFFRX1 f32_mux_0_data_reg_11_ ( .D(N433), .SI(f32_mux_0_data[10]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[11]) );
  SDFFRX1 f32_mux_0_data_reg_12_ ( .D(N434), .SI(f32_mux_0_data[11]), .SE(scan_enable), .CK(net121966), .RN(n859), .Q(f32_mux_0_data[12]) );
  SDFFRX1 f32_mux_0_data_reg_13_ ( .D(N435), .SI(f32_mux_0_data[12]), .SE(scan_enable), .CK(net121966), .RN(n860), .Q(f32_mux_0_data[13]) );
  SDFFRX1 f32_mux_0_data_reg_14_ ( .D(N436), .SI(f32_mux_0_data[13]), .SE(scan_enable), .CK(net121966), .RN(n861), .Q(f32_mux_0_data[14]) );
  SDFFRX1 f32_mux_0_data_reg_15_ ( .D(N437), .SI(f32_mux_0_data[14]), .SE(scan_enable), .CK(net121966), .RN(n129), .Q(f32_mux_0_data[15]) );
  SDFFX1 f32_data_reg_31_ ( .D(i_wr_data[31]), .SI(n_95_), .SE(scan_enable), .CK(net121977), .Q(n_94_) );
  SDFFX1 f32_data_reg_30_ ( .D(i_wr_data[30]), .SI(n_96_), .SE(scan_enable), .CK(net121977), .Q(n_95_) );
  SDFFX1 f32_data_reg_29_ ( .D(i_wr_data[29]), .SI(n_97_), .SE(scan_enable), .CK(net121977), .Q(n_96_) );
  SDFFX1 f32_data_reg_28_ ( .D(i_wr_data[28]), .SI(n_98_), .SE(scan_enable), .CK(net121977), .Q(n_97_) );
  SDFFX1 f32_data_reg_27_ ( .D(i_wr_data[27]), .SI(n_99_), .SE(scan_enable), .CK(net121977), .Q(n_98_) );
  SDFFX1 f32_data_reg_26_ ( .D(i_wr_data[26]), .SI(n_100_), .SE(scan_enable), .CK(net121977), .Q(n_99_) );
  SDFFX1 f32_data_reg_25_ ( .D(i_wr_data[25]), .SI(n_101_), .SE(scan_enable), .CK(net121977), .Q(n_100_) );
  SDFFX1 f32_data_reg_24_ ( .D(i_wr_data[24]), .SI(n_102_), .SE(scan_enable), .CK(net121977), .Q(n_101_) );
  SDFFX1 f32_data_reg_23_ ( .D(i_wr_data[23]), .SI(n_103_), .SE(scan_enable), .CK(net121977), .Q(n_102_) );
  SDFFX1 f32_data_reg_22_ ( .D(i_wr_data[22]), .SI(n_104_), .SE(scan_enable), .CK(net121977), .Q(n_103_) );
  SDFFX1 f32_data_reg_21_ ( .D(i_wr_data[21]), .SI(n_105_), .SE(scan_enable), .CK(net121977), .Q(n_104_) );
  SDFFX1 f32_data_reg_20_ ( .D(i_wr_data[20]), .SI(n_106_), .SE(scan_enable), .CK(net121977), .Q(n_105_) );
  SDFFX1 f32_data_reg_19_ ( .D(i_wr_data[19]), .SI(n_107_), .SE(scan_enable), .CK(net121977), .Q(n_106_) );
  SDFFX1 f32_data_reg_18_ ( .D(i_wr_data[18]), .SI(n_108_), .SE(scan_enable), .CK(net121977), .Q(n_107_) );
  SDFFX1 f32_data_reg_17_ ( .D(i_wr_data[17]), .SI(n_109_), .SE(scan_enable), .CK(net121977), .Q(n_108_) );
  SDFFX1 f32_data_reg_16_ ( .D(i_wr_data[16]), .SI(n_110_), .SE(scan_enable), .CK(net121977), .Q(n_109_) );
  SDFFX1 f32_data_reg_15_ ( .D(i_wr_data[15]), .SI(n_111_), .SE(scan_enable), .CK(net121977), .Q(n_110_) );
  SDFFX1 f32_data_reg_14_ ( .D(i_wr_data[14]), .SI(n_112_), .SE(scan_enable), .CK(net121977), .Q(n_111_) );
  SDFFX1 f32_data_reg_13_ ( .D(i_wr_data[13]), .SI(n_113_), .SE(scan_enable), .CK(net121977), .Q(n_112_) );
  SDFFX1 f32_data_reg_12_ ( .D(i_wr_data[12]), .SI(n_114_), .SE(scan_enable), .CK(net121977), .Q(n_113_) );
  SDFFX1 f32_data_reg_11_ ( .D(i_wr_data[11]), .SI(n1), .SE(scan_enable), .CK(net121977), .Q(n_114_) );
  SDFFX1 f32_data_reg_10_ ( .D(i_wr_data[10]), .SI(n_116_), .SE(scan_enable), .CK(net121977), .Q(test_so1) );
  SDFFX1 f32_data_reg_9_ ( .D(i_wr_data[9]), .SI(n_117_), .SE(scan_enable), .CK(net121977), .Q(n_116_) );
  SDFFX1 f32_data_reg_8_ ( .D(i_wr_data[8]), .SI(n_118_), .SE(scan_enable), .CK(net121977), .Q(n_117_) );
  SDFFX1 f32_data_reg_7_ ( .D(i_wr_data[7]), .SI(n_119_), .SE(scan_enable), .CK(net121977), .Q(n_118_) );
  SDFFX1 f32_data_reg_6_ ( .D(i_wr_data[6]), .SI(n_120_), .SE(scan_enable), .CK(net121977), .Q(n_119_) );
  SDFFX1 f32_data_reg_5_ ( .D(i_wr_data[5]), .SI(n_121_), .SE(scan_enable), .CK(net121977), .Q(n_120_) );
  SDFFX1 f32_data_reg_4_ ( .D(i_wr_data[4]), .SI(n_122_), .SE(scan_enable), .CK(net121977), .Q(n_121_) );
  SDFFX1 f32_data_reg_3_ ( .D(i_wr_data[3]), .SI(n_123_), .SE(scan_enable), .CK(net121977), .Q(n_122_) );
  SDFFX1 f32_data_reg_2_ ( .D(i_wr_data[2]), .SI(n_124_), .SE(scan_enable), .CK(net121977), .Q(n_123_) );
  SDFFX1 f32_data_reg_1_ ( .D(i_wr_data[1]), .SI(n_125_), .SE(scan_enable), .CK(net121977), .Q(n_124_) );
  SDFFX1 f32_data_reg_0_ ( .D(i_wr_data[0]), .SI(i_agg_su_count_a[31]), .SE(scan_enable), .CK(net121977), .Q(n_125_) );
  NOR2X2 U5 ( .A(n393), .B(n167), .Y(n836) );
  NOR2X2 U6 ( .A(n386), .B(n167), .Y(n843) );
  NOR3X4 U7 ( .A(n169), .B(n393), .C(n132), .Y(n857) );
  NOR3X2 U8 ( .A(n394), .B(n393), .C(n500), .Y(n674) );
  AND2X4 U9 ( .A(n845), .B(n852), .Y(n821) );
  NOR2X4 U10 ( .A(n380), .B(n383), .Y(n323) );
  NAND3X2 U11 ( .A(n370), .B(n369), .C(n371), .Y(n383) );
  INVX2 U15 ( .A(n126), .Y(n129) );
  INVX2 U16 ( .A(scan_iso_or2), .Y(n370) );
  BUFX8 U17 ( .A(n127), .Y(n861) );
  BUFX8 U18 ( .A(n127), .Y(n860) );
  BUFX8 U19 ( .A(n127), .Y(n859) );
  NAND3X2 U22 ( .A(n369), .B(scan_iso_or1), .C(scan_iso_or2), .Y(n167) );
  NAND3X2 U23 ( .A(n369), .B(n370), .C(scan_iso_or1), .Y(n160) );
  BUFX4 U24 ( .A(n674), .Y(n769) );
  NOR2X2 U26 ( .A(n393), .B(n373), .Y(n736) );
  BUFX4 U28 ( .A(n374), .Y(n130) );
  NOR2X4 U29 ( .A(o_reg_addr_reg_1__scan_iso_or_n), .B(o_reg_addr_reg_0__scan_iso_or_n), .Y(n131) );
  NAND3X2 U30 ( .A(scan_iso_or2), .B(scan_iso_or1), .C(n372), .Y(n373) );
  NOR2X2 U31 ( .A(n386), .B(n383), .Y(n374) );
  NOR2X1 U33 ( .A(n385), .B(n393), .Y(n839) );
  NOR2X4 U34 ( .A(scan_iso_or5), .B(n500), .Y(n852) );
  NOR2X1 U35 ( .A(n386), .B(n169), .Y(n845) );
  NOR2X1 U36 ( .A(n382), .B(n169), .Y(n846) );
  NOR2X1 U37 ( .A(n132), .B(n396), .Y(n823) );
  NOR2X1 U38 ( .A(n382), .B(n167), .Y(n831) );
  NOR2X1 U39 ( .A(n380), .B(n169), .Y(n847) );
  NOR2X1 U40 ( .A(n167), .B(n380), .Y(n844) );
  OR2X1 U41 ( .A(scan_iso_or4), .B(scan_iso_or3), .Y(n393) );
  NAND2X2 U42 ( .A(scan_iso_or5), .B(n131), .Y(n395) );
  OAI21X1 U44 ( .A0(n205), .A1(n204), .B0(n852), .Y(n209) );
  AND2X2 U45 ( .A(n846), .B(n852), .Y(n165) );
  OAI21X1 U46 ( .A0(n194), .A1(n193), .B0(n852), .Y(n198) );
  AND2X2 U47 ( .A(n831), .B(n852), .Y(n166) );
  AND2X2 U48 ( .A(n847), .B(n852), .Y(n170) );
  AND2X2 U49 ( .A(n844), .B(n852), .Y(n168) );
  NOR2X1 U50 ( .A(n132), .B(n210), .Y(n217) );
  BUFX4 U51 ( .A(n857), .Y(n814) );
  BUFX2 U52 ( .A(n821), .Y(n807) );
  AO22X1 U54 ( .A0(n769), .A1(i_hisbuf2_3[31]), .B0(n732), .B1(i_agg_su_count_a[31]), .Y(n504) );
  BUFX4 U55 ( .A(n492), .Y(n666) );
  AO22X1 U56 ( .A0(n769), .A1(i_hisbuf2_3[26]), .B0(n732), .B1(i_agg_su_count_a[26]), .Y(n488) );
  AO22X1 U57 ( .A0(n769), .A1(i_hisbuf2_3[25]), .B0(n732), .B1(i_agg_su_count_a[25]), .Y(n481) );
  AO22X1 U58 ( .A0(n769), .A1(i_hisbuf2_3[24]), .B0(n732), .B1(i_agg_su_count_a[24]), .Y(n496) );
  NOR2X1 U59 ( .A(n386), .B(n381), .Y(n710) );
  BUFX4 U60 ( .A(n711), .Y(n761) );
  BUFX4 U61 ( .A(n750), .Y(n656) );
  NOR2X2 U62 ( .A(scan_iso_or5), .B(n369), .Y(n372) );
  NOR2X1 U63 ( .A(n382), .B(n383), .Y(n829) );
  NOR2X2 U64 ( .A(scan_iso_or), .B(scan_iso_or1), .Y(n153) );
  NAND2X2 U65 ( .A(scan_iso_or3), .B(scan_iso_or4), .Y(n382) );
  NOR2X2 U66 ( .A(f_state[2]), .B(n152), .Y(n158) );
  INVX2 U67 ( .A(n323), .Y(n834) );
  NAND2X1 U68 ( .A(n852), .B(n158), .Y(n187) );
  NOR2X2 U69 ( .A(n335), .B(n_write), .Y(n336) );
  AO21X2 U70 ( .A0(n158), .A1(n157), .B0(f_err_ack), .Y(o_err_ack) );
  OAI31X1 U71 ( .A0(scan_iso_or5), .A1(n385), .A2(n386), .B0(n155), .Y(n157) );
  AOI21X1 U72 ( .A0(scan_iso_or5), .A1(n154), .B0(n500), .Y(n155) );
  OAI21X1 U73 ( .A0(n370), .A1(n382), .B0(n153), .Y(n154) );
  NAND2BX1 U75 ( .AN(f_state[1]), .B(f_state[0]), .Y(n152) );
  NOR2X1 U76 ( .A(n834), .B(n187), .Y(w_load_adj_config) );
  NOR2X1 U77 ( .A(n210), .B(n187), .Y(w_load_spare_config) );
  OAI21X1 U78 ( .A0(n230), .A1(n132), .B0(n229), .Y(N437) );
  OAI21X1 U79 ( .A0(n321), .A1(n132), .B0(n320), .Y(N436) );
  OAI21X1 U80 ( .A0(n310), .A1(n132), .B0(n309), .Y(N435) );
  OAI21X1 U81 ( .A0(n300), .A1(n132), .B0(n299), .Y(N434) );
  OAI21X1 U82 ( .A0(n240), .A1(n132), .B0(n239), .Y(N433) );
  OAI21X1 U83 ( .A0(n334), .A1(n132), .B0(n333), .Y(N432) );
  OAI21X1 U84 ( .A0(n260), .A1(n132), .B0(n259), .Y(N431) );
  OAI21X1 U85 ( .A0(n280), .A1(n132), .B0(n279), .Y(N430) );
  OAI21X1 U86 ( .A0(n250), .A1(n132), .B0(n249), .Y(N429) );
  OAI21X1 U87 ( .A0(n270), .A1(n132), .B0(n269), .Y(N428) );
  OAI21X1 U88 ( .A0(n290), .A1(n132), .B0(n289), .Y(N427) );
  OAI21X1 U89 ( .A0(n186), .A1(n132), .B0(n185), .Y(N426) );
  OAI21X1 U90 ( .A0(n176), .A1(n132), .B0(n175), .Y(N425) );
  NAND4X1 U91 ( .A(n209), .B(n208), .C(n207), .D(n206), .Y(N424) );
  NAND4X1 U92 ( .A(n198), .B(n197), .C(n196), .D(n195), .Y(N423) );
  NAND3X1 U93 ( .A(n828), .B(n827), .C(n826), .Y(N438) );
  NAND3X1 U94 ( .A(n348), .B(n347), .C(n346), .Y(N439) );
  NAND3X1 U95 ( .A(n792), .B(n791), .C(n790), .Y(N440) );
  AOI21X1 U96 ( .A0(n852), .A1(n789), .B0(n788), .Y(n790) );
  NAND3X1 U97 ( .A(n802), .B(n801), .C(n800), .Y(N441) );
  NAND3X1 U98 ( .A(n813), .B(n812), .C(n811), .Y(N442) );
  NAND3X1 U99 ( .A(n358), .B(n357), .C(n356), .Y(N443) );
  NAND3X1 U100 ( .A(n368), .B(n367), .C(n366), .Y(N444) );
  NAND3X1 U101 ( .A(n782), .B(n781), .C(n780), .Y(N445) );
  AOI21X1 U102 ( .A0(n852), .A1(n779), .B0(n778), .Y(n780) );
  NAND2X1 U103 ( .A(n212), .B(n211), .Y(N449) );
  NAND2X1 U104 ( .A(n220), .B(n219), .Y(N450) );
  NAND2X1 U105 ( .A(n216), .B(n215), .Y(N451) );
  NAND2X1 U106 ( .A(n214), .B(n213), .Y(N452) );
  NAND3X1 U107 ( .A(n507), .B(n506), .C(n505), .Y(N485) );
  NAND3X1 U108 ( .A(n454), .B(n453), .C(n452), .Y(N484) );
  NAND3X1 U109 ( .A(n473), .B(n472), .C(n471), .Y(N483) );
  NAND3X1 U110 ( .A(n470), .B(n469), .C(n468), .Y(N482) );
  NAND3X1 U111 ( .A(n477), .B(n476), .C(n475), .Y(N481) );
  NAND3X1 U112 ( .A(n491), .B(n490), .C(n489), .Y(N480) );
  NAND3X1 U113 ( .A(n484), .B(n483), .C(n482), .Y(N479) );
  NAND3X1 U114 ( .A(n499), .B(n498), .C(n497), .Y(N478) );
  NAND3X1 U115 ( .A(n399), .B(n398), .C(n397), .Y(N477) );
  NAND2X1 U116 ( .A(n656), .B(i_hisbuf2_4[23]), .Y(n399) );
  NAND3X1 U117 ( .A(n412), .B(n411), .C(n410), .Y(N476) );
  NAND2X1 U118 ( .A(n656), .B(i_hisbuf2_4[22]), .Y(n412) );
  NAND3X1 U119 ( .A(n559), .B(n558), .C(n557), .Y(N475) );
  NAND2X1 U120 ( .A(n750), .B(i_hisbuf2_4[21]), .Y(n559) );
  NAND3X1 U121 ( .A(n546), .B(n545), .C(n544), .Y(N474) );
  NAND2X1 U122 ( .A(n656), .B(i_hisbuf2_4[20]), .Y(n546) );
  NAND3X1 U123 ( .A(n520), .B(n519), .C(n518), .Y(N473) );
  NAND2X1 U124 ( .A(n656), .B(i_hisbuf2_4[19]), .Y(n520) );
  NAND3X1 U125 ( .A(n533), .B(n532), .C(n531), .Y(N472) );
  NAND2X1 U126 ( .A(n656), .B(i_hisbuf2_4[18]), .Y(n533) );
  NAND3X1 U127 ( .A(n573), .B(n572), .C(n571), .Y(N471) );
  NAND2X1 U128 ( .A(n656), .B(i_hisbuf2_4[17]), .Y(n573) );
  NAND3X1 U129 ( .A(n586), .B(n585), .C(n584), .Y(N470) );
  NAND2X1 U130 ( .A(n656), .B(i_hisbuf2_4[16]), .Y(n586) );
  NAND3X1 U131 ( .A(n600), .B(n599), .C(n598), .Y(N469) );
  NAND2X1 U132 ( .A(n750), .B(i_hisbuf2_4[15]), .Y(n600) );
  NAND3X1 U133 ( .A(n690), .B(n689), .C(n688), .Y(N468) );
  NAND2X1 U134 ( .A(n750), .B(i_hisbuf2_4[14]), .Y(n690) );
  NAND3X1 U135 ( .A(n749), .B(n748), .C(n747), .Y(N467) );
  NAND2X1 U136 ( .A(n750), .B(i_hisbuf2_4[13]), .Y(n749) );
  NAND3X1 U137 ( .A(n703), .B(n702), .C(n701), .Y(N466) );
  NAND2X1 U138 ( .A(n750), .B(i_hisbuf2_4[12]), .Y(n703) );
  NAND3X1 U139 ( .A(n735), .B(n734), .C(n733), .Y(N465) );
  NAND2X1 U140 ( .A(n750), .B(i_hisbuf2_4[11]), .Y(n735) );
  NAND3X1 U141 ( .A(n772), .B(n771), .C(n770), .Y(N464) );
  NAND2X1 U142 ( .A(n750), .B(i_hisbuf2_4[10]), .Y(n772) );
  NAND3X1 U143 ( .A(n720), .B(n719), .C(n718), .Y(N463) );
  NAND2X1 U144 ( .A(n750), .B(i_hisbuf2_4[9]), .Y(n720) );
  NAND3X1 U145 ( .A(n467), .B(n466), .C(n465), .Y(N462) );
  NAND2X1 U146 ( .A(n750), .B(i_hisbuf2_4[8]), .Y(n467) );
  NAND3X1 U147 ( .A(n438), .B(n437), .C(n436), .Y(N461) );
  NAND2X1 U148 ( .A(n750), .B(i_hisbuf2_4[7]), .Y(n438) );
  NAND3X1 U149 ( .A(n425), .B(n424), .C(n423), .Y(N460) );
  NAND2X1 U150 ( .A(n656), .B(i_hisbuf2_4[6]), .Y(n425) );
  NAND3X1 U151 ( .A(n626), .B(n625), .C(n624), .Y(N459) );
  NAND3X1 U152 ( .A(n677), .B(n676), .C(n675), .Y(N458) );
  NAND2X1 U153 ( .A(n656), .B(i_hisbuf2_4[4]), .Y(n677) );
  NAND3X1 U154 ( .A(n639), .B(n638), .C(n637), .Y(N457) );
  NAND2X1 U155 ( .A(n656), .B(i_hisbuf2_4[3]), .Y(n639) );
  NAND3X1 U156 ( .A(n655), .B(n654), .C(n653), .Y(N456) );
  NAND2X1 U157 ( .A(n656), .B(i_hisbuf2_4[2]), .Y(n655) );
  NAND3X1 U158 ( .A(n451), .B(n450), .C(n449), .Y(N455) );
  NAND3X1 U159 ( .A(n613), .B(n612), .C(n611), .Y(N454) );
  NAND2X1 U160 ( .A(n656), .B(i_hisbuf2_4[0]), .Y(n613) );
  NOR2X2 U161 ( .A(n385), .B(n380), .Y(n159) );
  NOR2X4 U162 ( .A(n380), .B(n373), .Y(n641) );
  AOI22X1 U163 ( .A0(n311), .A1(i_hisbuf0_1[2]), .B0(i_hisbuf3_1[2]), .B1(n843), .Y(n203) );
  AOI22X1 U164 ( .A0(n839), .A1(i_hb_sup[0]), .B0(n838), .B1(i_hisbuf1_0[0]), .Y(n840) );
  AOI22X1 U165 ( .A0(n815), .A1(i_hisbuf3_0[17]), .B0(n836), .B1(i_hisbuf2_1[17]), .Y(n340) );
  AOI22X1 U166 ( .A0(n815), .A1(i_hisbuf3_0[20]), .B0(n836), .B1(i_hisbuf2_1[20]), .Y(n805) );
  AOI22X1 U167 ( .A0(n311), .A1(i_hisbuf0_1[23]), .B0(n816), .B1(i_hisbuf1_1[23]), .Y(n774) );
  AOI22X1 U168 ( .A0(n751), .A1(i_hisbuf2_5[26]), .B0(i_hisbuf3_3[26]), .B1(n752), .Y(n486) );
  AOI22X1 U169 ( .A0(n640), .A1(i_hisbuf0_4[23]), .B0(n704), .B1(i_hisbuf3_3[23]), .Y(n377) );
  AOI22X1 U170 ( .A0(n753), .A1(i_hisbuf3_5[21]), .B0(n641), .B1(i_hisbuf0_6[21]), .Y(n548) );
  AOI22X1 U171 ( .A0(n642), .A1(i_hisbuf1_6[19]), .B0(n705), .B1(i_hisbuf3_6[19]), .Y(n508) );
  AOI22X1 U172 ( .A0(n663), .A1(i_hisbuf0_5[17]), .B0(n759), .B1(i_hisbuf3_4[17]), .Y(n568) );
  AOI22X1 U173 ( .A0(n564), .A1(i_hisbuf0_7[15]), .B0(n664), .B1(i_hisbuf1_5[15]), .Y(n593) );
  AOI22X1 U174 ( .A0(n666), .A1(i_hisbuf2_6[13]), .B0(n760), .B1(i_hisbuf2_7[13]), .Y(n742) );
  AOI22X1 U175 ( .A0(n667), .A1(i_hisbuf1_7[11]), .B0(n761), .B1(i_hisbuf3_7[11]), .Y(n725) );
  AOI22X1 U176 ( .A0(n657), .A1(i_hisbuf1_4[10]), .B0(n751), .B1(i_hisbuf2_5[10]), .Y(n758) );
  AOI22X1 U177 ( .A0(n640), .A1(i_hisbuf0_4[8]), .B0(n752), .B1(i_hisbuf3_3[8]), .Y(n457) );
  AOI22X1 U178 ( .A0(n642), .A1(i_hisbuf1_6[6]), .B0(n705), .B1(i_hisbuf3_6[6]), .Y(n413) );
  AOI22X1 U179 ( .A0(n564), .A1(i_hisbuf0_7[4]), .B0(n664), .B1(i_hisbuf1_5[4]), .Y(n670) );
  AOI22X1 U180 ( .A0(n640), .A1(i_hisbuf0_4[1]), .B0(n704), .B1(i_hisbuf3_3[1]), .Y(n441) );
  AOI22X1 U181 ( .A0(n311), .A1(i_hisbuf0_1[15]), .B0(n816), .B1(i_hisbuf1_1[15]), .Y(n222) );
  AOI22X1 U182 ( .A0(n165), .A1(i_hisbuf1_3[11]), .B0(n166), .B1(i_hisbuf1_2[11]), .Y(n238) );
  AOI22X1 U183 ( .A0(n168), .A1(i_hisbuf0_2[7]), .B0(n328), .B1(i_hisbuf3_1[7]), .Y(n246) );
  AOI22X1 U184 ( .A0(n170), .A1(i_hisbuf0_3[5]), .B0(i_hisbuf2_1[5]), .B1(n134), .Y(n285) );
  AOI22X1 U185 ( .A0(n838), .A1(i_hisbuf1_0[4]), .B0(i_hisbuf2_0[4]), .B1(n830), .Y(n180) );
  AO21X1 U186 ( .A0(n823), .A1(i_hisbuf0_0[21]), .B0(n353_inv), .Y(n354) );
  OA21X1 U187 ( .A0(f32_mux_0_data[4]), .A1(f32_mux_1_data[4]), .B0(n337), .Y(o_rd_data[4]) );
  OA21X1 U188 ( .A0(f32_mux_0_data[19]), .A1(f32_mux_1_data[19]), .B0(n337), .Y(o_rd_data[19]) );
  AOI22X1 U189 ( .A0(n168), .A1(i_hisbuf0_2[2]), .B0(n166), .B1(i_hisbuf1_2[2]), .Y(n207) );
  AOI22X1 U190 ( .A0(n814), .A1(i_hisbuf2_2[28]), .B0(i_hisbuf2_1[28]), .B1(n134), .Y(n220) );
  AOI22X1 U191 ( .A0(n732), .A1(i_agg_su_count_a[29]), .B0(n760), .B1(i_hisbuf2_7[29]), .Y(n471) );
  AOI22X1 U192 ( .A0(n769), .A1(i_hisbuf2_3[19]), .B0(n768), .B1(i_agg_su_count_a[19]), .Y(n518) );
  AOI22X1 U193 ( .A0(n769), .A1(i_hisbuf2_3[14]), .B0(n732), .B1(i_agg_su_count_a[14]), .Y(n688) );
  AOI22X1 U194 ( .A0(n769), .A1(i_hisbuf2_3[9]), .B0(n768), .B1(i_agg_su_count_a[9]), .Y(n718) );
  INVX2 U195 ( .A(scan_iso_or), .Y(n369) );
  INVX2 U196 ( .A(scan_iso_or1), .Y(n371) );
  NOR2X2 U197 ( .A(n386), .B(n160), .Y(n837) );
  NOR2X2 U198 ( .A(n393), .B(n160), .Y(n322) );
  BUFX4 U199 ( .A(n322), .Y(n830) );
  AO22X1 U200 ( .A0(n837), .A1(i_hisbuf3_0[27]), .B0(n830), .B1(i_hisbuf2_0[31]), .Y(n133) );
  AOI21X1 U201 ( .A0(n374), .A1(i_spare_config[31]), .B0(n133), .Y(n137) );
  AOI22X1 U203 ( .A0(n807), .A1(i_hisbuf3_2[27]), .B0(i_hisbuf2_1[31]), .B1(n134), .Y(n136) );
  AOI22X1 U205 ( .A0(n857), .A1(i_hisbuf2_2[31]), .B0(n328), .B1(i_hisbuf3_1[27]), .Y(n135) );
  OAI211X1 U206 ( .A0(n132), .A1(n137), .B0(n136), .C0(n135), .Y(N453) );
  AO22X1 U208 ( .A0(n815), .A1(i_hisbuf3_0[24]), .B0(n830), .B1(i_hisbuf2_0[24]), .Y(n138) );
  AOI21X1 U209 ( .A0(n374), .A1(i_spare_config[24]), .B0(n138), .Y(n141) );
  AOI22X1 U210 ( .A0(n807), .A1(i_hisbuf3_2[24]), .B0(i_hisbuf2_1[24]), .B1(n134), .Y(n140) );
  AOI22X1 U211 ( .A0(n857), .A1(i_hisbuf2_2[24]), .B0(n328), .B1(i_hisbuf3_1[24]), .Y(n139) );
  OAI211X1 U212 ( .A0(n132), .A1(n141), .B0(n140), .C0(n139), .Y(N446) );
  AO22X1 U213 ( .A0(n815), .A1(i_hisbuf3_0[26]), .B0(n830), .B1(i_hisbuf2_0[26]), .Y(n142) );
  AOI21X1 U214 ( .A0(n374), .A1(i_spare_config[26]), .B0(n142), .Y(n145) );
  AOI22X1 U215 ( .A0(n807), .A1(i_hisbuf3_2[26]), .B0(i_hisbuf2_1[26]), .B1(n134), .Y(n144) );
  AOI22X1 U216 ( .A0(n857), .A1(i_hisbuf2_2[26]), .B0(n328), .B1(i_hisbuf3_1[26]), .Y(n143) );
  OAI211X1 U217 ( .A0(n132), .A1(n145), .B0(n144), .C0(n143), .Y(N448) );
  AO22X1 U218 ( .A0(n815), .A1(i_hisbuf3_0[25]), .B0(n830), .B1(i_hisbuf2_0[25]), .Y(n146) );
  AOI21X1 U219 ( .A0(n374), .A1(i_spare_config[25]), .B0(n146), .Y(n149) );
  AOI22X1 U220 ( .A0(n807), .A1(i_hisbuf3_2[25]), .B0(i_hisbuf2_1[25]), .B1(n134), .Y(n148) );
  AOI22X1 U221 ( .A0(n857), .A1(i_hisbuf2_2[25]), .B0(n328), .B1(i_hisbuf3_1[25]), .Y(n147) );
  OAI211X1 U222 ( .A0(n132), .A1(n149), .B0(n148), .C0(n147), .Y(N447) );
  NOR2X1 U223 ( .A(i_rd_strb), .B(i_wr_strb), .Y(n150) );
  NAND2X1 U224 ( .A(n152), .B(n150), .Y(N405) );
  INVX2 U225 ( .A(n150), .Y(N410) );
  NOR2X1 U226 ( .A(n152), .B(N410), .Y(N406) );
  NAND2BX1 U227 ( .AN(n152), .B(f_state[2]), .Y(n156) );
  INVX2 U228 ( .A(i_rd_strb), .Y(n151) );
  AOI21X1 U229 ( .A0(n156), .A1(n151), .B0(i_wr_strb), .Y(N407) );
  NOR2X1 U230 ( .A(n156), .B(N410), .Y(N408) );
  AO21X1 U231 ( .A0(n_write), .A1(n335), .B0(i_wr_strb), .Y(n842) );
  NAND2X4 U232 ( .A(scan_iso_or2), .B(n153), .Y(n385) );
  NOR2X1 U233 ( .A(n157), .B(n156), .Y(N420) );
  INVX2 U234 ( .A(n156), .Y(N421) );
  AND2X1 U235 ( .A(n157), .B(N421), .Y(N409) );
  INVX2 U236 ( .A(n829), .Y(n384) );
  NOR2X1 U237 ( .A(n384), .B(n187), .Y(w_load_dbg_config) );
  INVX2 U238 ( .A(n374), .Y(n210) );
  INVX2 U239 ( .A(n335), .Y(o_ack) );
  NOR2X4 U240 ( .A(n385), .B(n382), .Y(n838) );
  AOI22X1 U241 ( .A0(n838), .A1(i_hisbuf1_0[3]), .B0(i_hisbuf2_0[3]), .B1(n830), .Y(n164) );
  NAND2BX4 U242 ( .AN(scan_iso_or4), .B(scan_iso_or3), .Y(n380) );
  AOI22X1 U243 ( .A0(n837), .A1(i_hisbuf3_0[3]), .B0(n159), .B1(i_hisbuf0_0[3]), .Y(n163) );
  NOR2X4 U244 ( .A(n160), .B(n380), .Y(n311) );
  NOR2X4 U245 ( .A(n382), .B(n160), .Y(n816) );
  AOI22X1 U246 ( .A0(n311), .A1(i_hisbuf0_1[3]), .B0(n816), .B1(i_hisbuf1_1[3]), .Y(n162) );
  AOI22X1 U247 ( .A0(n323), .A1(scan_iso_or9), .B0(n130), .B1(i_spare_config[3]), .Y(n161) );
  AND4X1 U248 ( .A(n164), .B(n163), .C(n162), .D(n161), .Y(n176) );
  AOI22X1 U249 ( .A0(n165), .A1(i_hisbuf1_3[3]), .B0(n166), .B1(i_hisbuf1_2[3]), .Y(n174) );
  AOI22X1 U250 ( .A0(n857), .A1(i_hisbuf2_2[3]), .B0(n821), .B1(i_hisbuf3_2[3]), .Y(n173) );
  AOI22X1 U251 ( .A0(n168), .A1(i_hisbuf0_2[3]), .B0(n328), .B1(i_hisbuf3_1[3]), .Y(n172) );
  AOI22X1 U252 ( .A0(n170), .A1(i_hisbuf0_3[3]), .B0(i_hisbuf2_1[3]), .B1(n134), .Y(n171) );
  AND4X1 U253 ( .A(n174), .B(n173), .C(n172), .D(n171), .Y(n175) );
  AOI22X1 U254 ( .A0(n837), .A1(i_hisbuf3_0[4]), .B0(n159), .B1(i_hisbuf0_0[4]), .Y(n179) );
  AOI22X1 U255 ( .A0(n311), .A1(i_hisbuf0_1[4]), .B0(n816), .B1(i_hisbuf1_1[4]), .Y(n178) );
  AOI22X1 U256 ( .A0(n323), .A1(o_adj_config[4]), .B0(n130), .B1(i_spare_config[4]), .Y(n177) );
  AND4X1 U257 ( .A(n180), .B(n179), .C(n178), .D(n177), .Y(n186) );
  AOI22X1 U258 ( .A0(n165), .A1(i_hisbuf1_3[4]), .B0(n166), .B1(i_hisbuf1_2[4]), .Y(n184) );
  AOI22X1 U259 ( .A0(n857), .A1(i_hisbuf2_2[4]), .B0(n807), .B1(i_hisbuf3_2[4]), .Y(n183) );
  AOI22X1 U260 ( .A0(n168), .A1(i_hisbuf0_2[4]), .B0(n328), .B1(i_hisbuf3_1[4]), .Y(n182) );
  AOI22X1 U261 ( .A0(n170), .A1(i_hisbuf0_3[4]), .B0(i_hisbuf2_1[4]), .B1(n134), .Y(n181) );
  AND4X1 U262 ( .A(n184), .B(n183), .C(n182), .D(n181), .Y(n185) );
  AOI22X1 U263 ( .A0(n839), .A1(i_hb_sup[1]), .B0(n130), .B1(i_spare_config[1]), .Y(n188) );
  AO21X1 U264 ( .A0(n838), .A1(i_hisbuf1_0[1]), .B0(n188_inv), .Y(n194) );
  AOI22X1 U265 ( .A0(n311), .A1(i_hisbuf0_1[1]), .B0(i_hisbuf3_1[1]), .B1(n843), .Y(n192) );
  AOI22X1 U266 ( .A0(n816), .A1(i_hisbuf1_1[1]), .B0(n323), .B1(scan_iso_or6), .Y(n191) );
  AOI22X1 U267 ( .A0(n815), .A1(i_hisbuf3_0[1]), .B0(n159), .B1(i_hisbuf0_0[1]), .Y(n190) );
  AOI22X1 U268 ( .A0(n836), .A1(i_hisbuf2_1[1]), .B0(i_hisbuf2_0[1]), .B1(n830), .Y(n189) );
  NAND4X1 U269 ( .A(n192), .B(n191), .C(n190), .D(n189), .Y(n193) );
  AOI22X1 U270 ( .A0(n170), .A1(i_hisbuf0_3[1]), .B0(n165), .B1(i_hisbuf1_3[1]), .Y(n197) );
  AOI22X1 U271 ( .A0(n168), .A1(i_hisbuf0_2[1]), .B0(n166), .B1(i_hisbuf1_2[1]), .Y(n196) );
  AOI22X1 U272 ( .A0(n814), .A1(i_hisbuf2_2[1]), .B0(n821), .B1(i_hisbuf3_2[1]), .Y(n195) );
  AOI22X1 U273 ( .A0(n839), .A1(i_hb_sup[2]), .B0(n130), .B1(i_spare_config[2]), .Y(n199) );
  AO21X1 U274 ( .A0(n838), .A1(i_hisbuf1_0[2]), .B0(n199_inv), .Y(n205) );
  AOI22X1 U275 ( .A0(n816), .A1(i_hisbuf1_1[2]), .B0(n323), .B1(scan_iso_or8), .Y(n202) );
  AOI22X1 U276 ( .A0(n815), .A1(i_hisbuf3_0[2]), .B0(n159), .B1(i_hisbuf0_0[2]), .Y(n201) );
  AOI22X1 U277 ( .A0(n836), .A1(i_hisbuf2_1[2]), .B0(i_hisbuf2_0[2]), .B1(n830), .Y(n200) );
  NAND4X1 U278 ( .A(n203), .B(n202), .C(n201), .D(n200), .Y(n204) );
  AOI22X1 U279 ( .A0(n170), .A1(i_hisbuf0_3[2]), .B0(n165), .B1(i_hisbuf1_3[2]), .Y(n208) );
  AOI22X1 U280 ( .A0(n814), .A1(i_hisbuf2_2[2]), .B0(n821), .B1(i_hisbuf3_2[2]), .Y(n206) );
  AOI22X1 U281 ( .A0(n814), .A1(i_hisbuf2_2[27]), .B0(i_hisbuf2_1[27]), .B1(n134), .Y(n212) );
  AND2X1 U282 ( .B(n830), .A(n132_inv), .Y(n218) );
  INVX1 U282_inv ( .A(n132), .Y(n132_inv) );
  AOI22X1 U283 ( .A0(n218), .A1(i_hisbuf2_0[27]), .B0(n217), .B1(i_spare_config[27]), .Y(n211) );
  AOI22X1 U284 ( .A0(n814), .A1(i_hisbuf2_2[30]), .B0(i_hisbuf2_1[30]), .B1(n134), .Y(n214) );
  AOI22X1 U285 ( .A0(n218), .A1(i_hisbuf2_0[30]), .B0(n217), .B1(i_spare_config[30]), .Y(n213) );
  AOI22X1 U286 ( .A0(n814), .A1(i_hisbuf2_2[29]), .B0(i_hisbuf2_1[29]), .B1(n134), .Y(n216) );
  AOI22X1 U287 ( .A0(n218), .A1(i_hisbuf2_0[29]), .B0(n217), .B1(i_spare_config[29]), .Y(n215) );
  AOI22X1 U288 ( .A0(n218), .A1(i_hisbuf2_0[28]), .B0(n217), .B1(i_spare_config[28]), .Y(n219) );
  AOI22X1 U289 ( .A0(n838), .A1(i_hisbuf1_0[15]), .B0(i_hisbuf2_0[15]), .B1(n322), .Y(n224) );
  AOI22X1 U290 ( .A0(n815), .A1(i_hisbuf3_0[15]), .B0(n159), .B1(i_hisbuf0_0[15]), .Y(n223) );
  AOI22X1 U291 ( .A0(n323), .A1(o_adj_config[15]), .B0(n130), .B1(i_spare_config[15]), .Y(n221) );
  AND4X1 U292 ( .A(n224), .B(n223), .C(n222), .D(n221), .Y(n230) );
  AOI22X1 U293 ( .A0(n165), .A1(i_hisbuf1_3[15]), .B0(n166), .B1(i_hisbuf1_2[15]), .Y(n228) );
  AOI22X1 U294 ( .A0(n814), .A1(i_hisbuf2_2[15]), .B0(n821), .B1(i_hisbuf3_2[15]), .Y(n227) );
  AOI22X1 U295 ( .A0(n168), .A1(i_hisbuf0_2[15]), .B0(n328), .B1(i_hisbuf3_1[15]), .Y(n226) );
  AOI22X1 U296 ( .A0(n170), .A1(i_hisbuf0_3[15]), .B0(i_hisbuf2_1[15]), .B1(n134), .Y(n225) );
  AND4X1 U297 ( .A(n228), .B(n227), .C(n226), .D(n225), .Y(n229) );
  AOI22X1 U298 ( .A0(n838), .A1(i_hisbuf1_0[11]), .B0(i_hisbuf2_0[11]), .B1(n322), .Y(n234) );
  AOI22X1 U299 ( .A0(n815), .A1(i_hisbuf3_0[11]), .B0(n159), .B1(i_hisbuf0_0[11]), .Y(n233) );
  AOI22X1 U300 ( .A0(n311), .A1(i_hisbuf0_1[11]), .B0(n816), .B1(i_hisbuf1_1[11]), .Y(n232) );
  AOI22X1 U301 ( .A0(n323), .A1(o_adj_config[11]), .B0(n130), .B1(i_spare_config[11]), .Y(n231) );
  AND4X1 U302 ( .A(n234), .B(n233), .C(n232), .D(n231), .Y(n240) );
  AOI22X1 U303 ( .A0(n814), .A1(i_hisbuf2_2[11]), .B0(n821), .B1(i_hisbuf3_2[11]), .Y(n237) );
  AOI22X1 U304 ( .A0(n168), .A1(i_hisbuf0_2[11]), .B0(n328), .B1(i_hisbuf3_1[11]), .Y(n236) );
  AOI22X1 U305 ( .A0(n170), .A1(i_hisbuf0_3[11]), .B0(i_hisbuf2_1[11]), .B1(n134), .Y(n235) );
  AND4X1 U306 ( .A(n238), .B(n237), .C(n236), .D(n235), .Y(n239) );
  AOI22X1 U307 ( .A0(n838), .A1(i_hisbuf1_0[7]), .B0(i_hisbuf2_0[7]), .B1(n830), .Y(n244) );
  AOI22X1 U308 ( .A0(n837), .A1(i_hisbuf3_0[7]), .B0(n159), .B1(i_hisbuf0_0[7]), .Y(n243) );
  AOI22X1 U309 ( .A0(n311), .A1(i_hisbuf0_1[7]), .B0(n816), .B1(i_hisbuf1_1[7]), .Y(n242) );
  AOI22X1 U310 ( .A0(n323), .A1(o_adj_config[7]), .B0(n130), .B1(i_spare_config[7]), .Y(n241) );
  AND4X1 U311 ( .A(n244), .B(n243), .C(n242), .D(n241), .Y(n250) );
  AOI22X1 U312 ( .A0(n165), .A1(i_hisbuf1_3[7]), .B0(n166), .B1(i_hisbuf1_2[7]), .Y(n248) );
  AOI22X1 U313 ( .A0(n814), .A1(i_hisbuf2_2[7]), .B0(n821), .B1(i_hisbuf3_2[7]), .Y(n247) );
  AOI22X1 U314 ( .A0(n170), .A1(i_hisbuf0_3[7]), .B0(i_hisbuf2_1[7]), .B1(n134), .Y(n245) );
  AND4X1 U315 ( .A(n248), .B(n247), .C(n246), .D(n245), .Y(n249) );
  AOI22X1 U316 ( .A0(n838), .A1(i_hisbuf1_0[9]), .B0(i_hisbuf2_0[9]), .B1(n830), .Y(n254) );
  AOI22X1 U317 ( .A0(n815), .A1(i_hisbuf3_0[9]), .B0(n159), .B1(i_hisbuf0_0[9]), .Y(n253) );
  AOI22X1 U318 ( .A0(n311), .A1(i_hisbuf0_1[9]), .B0(n816), .B1(i_hisbuf1_1[9]), .Y(n252) );
  AOI22X1 U319 ( .A0(n323), .A1(o_adj_config[9]), .B0(n130), .B1(i_spare_config[9]), .Y(n251) );
  AND4X1 U320 ( .A(n254), .B(n253), .C(n252), .D(n251), .Y(n260) );
  AOI22X1 U321 ( .A0(n165), .A1(i_hisbuf1_3[9]), .B0(n166), .B1(i_hisbuf1_2[9]), .Y(n258) );
  AOI22X1 U322 ( .A0(n814), .A1(i_hisbuf2_2[9]), .B0(n821), .B1(i_hisbuf3_2[9]), .Y(n257) );
  AOI22X1 U323 ( .A0(n168), .A1(i_hisbuf0_2[9]), .B0(n328), .B1(i_hisbuf3_1[9]), .Y(n256) );
  AOI22X1 U324 ( .A0(n170), .A1(i_hisbuf0_3[9]), .B0(i_hisbuf2_1[9]), .B1(n134), .Y(n255) );
  AND4X1 U325 ( .A(n258), .B(n257), .C(n256), .D(n255), .Y(n259) );
  AOI22X1 U326 ( .A0(n838), .A1(i_hisbuf1_0[6]), .B0(i_hisbuf2_0[6]), .B1(n322), .Y(n264) );
  AOI22X1 U327 ( .A0(n837), .A1(i_hisbuf3_0[6]), .B0(n159), .B1(i_hisbuf0_0[6]), .Y(n263) );
  AOI22X1 U328 ( .A0(n311), .A1(i_hisbuf0_1[6]), .B0(n816), .B1(i_hisbuf1_1[6]), .Y(n262) );
  AOI22X1 U329 ( .A0(n323), .A1(o_adj_config[6]), .B0(n130), .B1(i_spare_config[6]), .Y(n261) );
  AND4X1 U330 ( .A(n264), .B(n263), .C(n262), .D(n261), .Y(n270) );
  AOI22X1 U331 ( .A0(n165), .A1(i_hisbuf1_3[6]), .B0(n166), .B1(i_hisbuf1_2[6]), .Y(n268) );
  AOI22X1 U332 ( .A0(n814), .A1(i_hisbuf2_2[6]), .B0(n821), .B1(i_hisbuf3_2[6]), .Y(n267) );
  AOI22X1 U333 ( .A0(n168), .A1(i_hisbuf0_2[6]), .B0(n328), .B1(i_hisbuf3_1[6]), .Y(n266) );
  AOI22X1 U334 ( .A0(n170), .A1(i_hisbuf0_3[6]), .B0(i_hisbuf2_1[6]), .B1(n134), .Y(n265) );
  AND4X1 U335 ( .A(n268), .B(n267), .C(n266), .D(n265), .Y(n269) );
  AOI22X1 U336 ( .A0(n838), .A1(i_hisbuf1_0[8]), .B0(i_hisbuf2_0[8]), .B1(n830), .Y(n274) );
  AOI22X1 U337 ( .A0(n815), .A1(i_hisbuf3_0[8]), .B0(n159), .B1(i_hisbuf0_0[8]), .Y(n273) );
  AOI22X1 U338 ( .A0(n311), .A1(i_hisbuf0_1[8]), .B0(n816), .B1(i_hisbuf1_1[8]), .Y(n272) );
  AOI22X1 U339 ( .A0(n323), .A1(o_adj_config[8]), .B0(n130), .B1(i_spare_config[8]), .Y(n271) );
  AND4X1 U340 ( .A(n274), .B(n273), .C(n272), .D(n271), .Y(n280) );
  AOI22X1 U341 ( .A0(n165), .A1(i_hisbuf1_3[8]), .B0(n166), .B1(i_hisbuf1_2[8]), .Y(n278) );
  AOI22X1 U342 ( .A0(n814), .A1(i_hisbuf2_2[8]), .B0(n821), .B1(i_hisbuf3_2[8]), .Y(n277) );
  AOI22X1 U343 ( .A0(n168), .A1(i_hisbuf0_2[8]), .B0(n328), .B1(i_hisbuf3_1[8]), .Y(n276) );
  AOI22X1 U344 ( .A0(n170), .A1(i_hisbuf0_3[8]), .B0(i_hisbuf2_1[8]), .B1(n134), .Y(n275) );
  AND4X1 U345 ( .A(n278), .B(n277), .C(n276), .D(n275), .Y(n279) );
  AOI22X1 U346 ( .A0(n838), .A1(i_hisbuf1_0[5]), .B0(i_hisbuf2_0[5]), .B1(n830), .Y(n284) );
  AOI22X1 U347 ( .A0(n837), .A1(i_hisbuf3_0[5]), .B0(n159), .B1(i_hisbuf0_0[5]), .Y(n283) );
  AOI22X1 U348 ( .A0(n311), .A1(i_hisbuf0_1[5]), .B0(n816), .B1(i_hisbuf1_1[5]), .Y(n282) );
  AOI22X1 U349 ( .A0(n323), .A1(o_adj_config[5]), .B0(n130), .B1(i_spare_config[5]), .Y(n281) );
  AND4X1 U350 ( .A(n284), .B(n283), .C(n282), .D(n281), .Y(n290) );
  AOI22X1 U351 ( .A0(n165), .A1(i_hisbuf1_3[5]), .B0(n166), .B1(i_hisbuf1_2[5]), .Y(n288) );
  AOI22X1 U352 ( .A0(n814), .A1(i_hisbuf2_2[5]), .B0(n821), .B1(i_hisbuf3_2[5]), .Y(n287) );
  AOI22X1 U353 ( .A0(n168), .A1(i_hisbuf0_2[5]), .B0(n328), .B1(i_hisbuf3_1[5]), .Y(n286) );
  AND4X1 U354 ( .A(n288), .B(n287), .C(n286), .D(n285), .Y(n289) );
  AOI22X1 U355 ( .A0(n838), .A1(i_hisbuf1_0[12]), .B0(i_hisbuf2_0[12]), .B1(n322), .Y(n294) );
  AOI22X1 U356 ( .A0(n815), .A1(i_hisbuf3_0[12]), .B0(n159), .B1(i_hisbuf0_0[12]), .Y(n293) );
  AOI22X1 U357 ( .A0(n311), .A1(i_hisbuf0_1[12]), .B0(n816), .B1(i_hisbuf1_1[12]), .Y(n292) );
  AOI22X1 U358 ( .A0(n323), .A1(o_adj_config[12]), .B0(n130), .B1(i_spare_config[12]), .Y(n291) );
  AND4X1 U359 ( .A(n294), .B(n293), .C(n292), .D(n291), .Y(n300) );
  AOI22X1 U360 ( .A0(n165), .A1(i_hisbuf1_3[12]), .B0(n166), .B1(i_hisbuf1_2[12]), .Y(n298) );
  AOI22X1 U361 ( .A0(n814), .A1(i_hisbuf2_2[12]), .B0(n821), .B1(i_hisbuf3_2[12]), .Y(n297) );
  AOI22X1 U362 ( .A0(n168), .A1(i_hisbuf0_2[12]), .B0(n328), .B1(i_hisbuf3_1[12]), .Y(n296) );
  AOI22X1 U363 ( .A0(n170), .A1(i_hisbuf0_3[12]), .B0(i_hisbuf2_1[12]), .B1(n134), .Y(n295) );
  AND4X1 U364 ( .A(n298), .B(n297), .C(n296), .D(n295), .Y(n299) );
  AOI22X1 U365 ( .A0(n838), .A1(i_hisbuf1_0[13]), .B0(i_hisbuf2_0[13]), .B1(n322), .Y(n304) );
  AOI22X1 U366 ( .A0(n815), .A1(i_hisbuf3_0[13]), .B0(n159), .B1(i_hisbuf0_0[13]), .Y(n303) );
  AOI22X1 U367 ( .A0(n311), .A1(i_hisbuf0_1[13]), .B0(n816), .B1(i_hisbuf1_1[13]), .Y(n302) );
  AOI22X1 U368 ( .A0(n323), .A1(o_adj_config[13]), .B0(n130), .B1(i_spare_config[13]), .Y(n301) );
  AND4X1 U369 ( .A(n304), .B(n303), .C(n302), .D(n301), .Y(n310) );
  AOI22X1 U370 ( .A0(n165), .A1(i_hisbuf1_3[13]), .B0(n166), .B1(i_hisbuf1_2[13]), .Y(n308) );
  AOI22X1 U371 ( .A0(n814), .A1(i_hisbuf2_2[13]), .B0(n821), .B1(i_hisbuf3_2[13]), .Y(n307) );
  AOI22X1 U372 ( .A0(n168), .A1(i_hisbuf0_2[13]), .B0(n328), .B1(i_hisbuf3_1[13]), .Y(n306) );
  AOI22X1 U373 ( .A0(n170), .A1(i_hisbuf0_3[13]), .B0(i_hisbuf2_1[13]), .B1(n134), .Y(n305) );
  AND4X1 U374 ( .A(n308), .B(n307), .C(n306), .D(n305), .Y(n309) );
  AOI22X1 U375 ( .A0(n838), .A1(i_hisbuf1_0[14]), .B0(i_hisbuf2_0[14]), .B1(n322), .Y(n315) );
  AOI22X1 U376 ( .A0(n815), .A1(i_hisbuf3_0[14]), .B0(n159), .B1(i_hisbuf0_0[14]), .Y(n314) );
  AOI22X1 U377 ( .A0(n311), .A1(i_hisbuf0_1[14]), .B0(n816), .B1(i_hisbuf1_1[14]), .Y(n313) );
  AOI22X1 U378 ( .A0(n323), .A1(o_adj_config[14]), .B0(n130), .B1(i_spare_config[14]), .Y(n312) );
  AND4X1 U379 ( .A(n315), .B(n314), .C(n313), .D(n312), .Y(n321) );
  AOI22X1 U380 ( .A0(n165), .A1(i_hisbuf1_3[14]), .B0(n166), .B1(i_hisbuf1_2[14]), .Y(n319) );
  AOI22X1 U381 ( .A0(n814), .A1(i_hisbuf2_2[14]), .B0(n821), .B1(i_hisbuf3_2[14]), .Y(n318) );
  AOI22X1 U382 ( .A0(n168), .A1(i_hisbuf0_2[14]), .B0(n328), .B1(i_hisbuf3_1[14]), .Y(n317) );
  AOI22X1 U383 ( .A0(n170), .A1(i_hisbuf0_3[14]), .B0(i_hisbuf2_1[14]), .B1(n134), .Y(n316) );
  AND4X1 U384 ( .A(n319), .B(n318), .C(n317), .D(n316), .Y(n320) );
  AOI22X1 U385 ( .A0(n838), .A1(i_hisbuf1_0[10]), .B0(i_hisbuf2_0[10]), .B1(n322), .Y(n327) );
  AOI22X1 U386 ( .A0(n815), .A1(i_hisbuf3_0[10]), .B0(n159), .B1(i_hisbuf0_0[10]), .Y(n326) );
  AOI22X1 U387 ( .A0(n311), .A1(i_hisbuf0_1[10]), .B0(n816), .B1(i_hisbuf1_1[10]), .Y(n325) );
  AOI22X1 U388 ( .A0(n323), .A1(o_adj_config[10]), .B0(n130), .B1(i_spare_config[10]), .Y(n324) );
  AND4X1 U389 ( .A(n327), .B(n326), .C(n325), .D(n324), .Y(n334) );
  AOI22X1 U390 ( .A0(n165), .A1(i_hisbuf1_3[10]), .B0(n166), .B1(i_hisbuf1_2[10]), .Y(n332) );
  AOI22X1 U391 ( .A0(n814), .A1(i_hisbuf2_2[10]), .B0(n821), .B1(i_hisbuf3_2[10]), .Y(n331) );
  AOI22X1 U392 ( .A0(n168), .A1(i_hisbuf0_2[10]), .B0(n328), .B1(i_hisbuf3_1[10]), .Y(n330) );
  AOI22X1 U393 ( .A0(n170), .A1(i_hisbuf0_3[10]), .B0(i_hisbuf2_1[10]), .B1(n134), .Y(n329) );
  AND4X1 U394 ( .A(n332), .B(n331), .C(n330), .D(n329), .Y(n333) );
  BUFX4 U395 ( .A(n336), .Y(n337) );
  OA21X1 U396 ( .A0(f32_mux_0_data[18]), .A1(f32_mux_1_data[18]), .B0(n337), .Y(o_rd_data[18]) );
  OA21X1 U397 ( .A0(f32_mux_0_data[21]), .A1(f32_mux_1_data[21]), .B0(n337), .Y(o_rd_data[21]) );
  OA21X1 U398 ( .A0(f32_mux_0_data[22]), .A1(f32_mux_1_data[22]), .B0(n337), .Y(o_rd_data[22]) );
  OA21X1 U399 ( .A0(f32_mux_0_data[20]), .A1(f32_mux_1_data[20]), .B0(n337), .Y(o_rd_data[20]) );
  OA21X1 U400 ( .A0(f32_mux_0_data[24]), .A1(f32_mux_1_data[24]), .B0(n336), .Y(o_rd_data[24]) );
  OA21X1 U401 ( .A0(f32_mux_0_data[23]), .A1(f32_mux_1_data[23]), .B0(n337), .Y(o_rd_data[23]) );
  OA21X1 U402 ( .A0(f32_mux_0_data[14]), .A1(f32_mux_1_data[14]), .B0(n337), .Y(o_rd_data[14]) );
  OA21X1 U403 ( .A0(f32_mux_0_data[25]), .A1(f32_mux_1_data[25]), .B0(n336), .Y(o_rd_data[25]) );
  OA21X1 U404 ( .A0(f32_mux_0_data[28]), .A1(f32_mux_1_data[28]), .B0(n337), .Y(o_rd_data[28]) );
  OA21X1 U405 ( .A0(f32_mux_0_data[26]), .A1(f32_mux_1_data[26]), .B0(n337), .Y(o_rd_data[26]) );
  OA21X1 U406 ( .A0(f32_mux_0_data[29]), .A1(f32_mux_1_data[29]), .B0(n336), .Y(o_rd_data[29]) );
  OA21X1 U407 ( .A0(f32_mux_0_data[27]), .A1(f32_mux_1_data[27]), .B0(n337), .Y(o_rd_data[27]) );
  OA21X1 U408 ( .A0(f32_mux_0_data[3]), .A1(f32_mux_1_data[3]), .B0(n337), .Y(o_rd_data[3]) );
  OA21X1 U409 ( .A0(f32_mux_0_data[2]), .A1(f32_mux_1_data[2]), .B0(n337), .Y(o_rd_data[2]) );
  OA21X1 U410 ( .A0(f32_mux_0_data[0]), .A1(f32_mux_1_data[0]), .B0(n337), .Y(o_rd_data[0]) );
  OA21X1 U411 ( .A0(f32_mux_0_data[30]), .A1(f32_mux_1_data[30]), .B0(n336), .Y(o_rd_data[30]) );
  OA21X1 U412 ( .A0(f32_mux_0_data[16]), .A1(f32_mux_1_data[16]), .B0(n336), .Y(o_rd_data[16]) );
  OA21X1 U413 ( .A0(f32_mux_0_data[31]), .A1(f32_mux_1_data[31]), .B0(n336), .Y(o_rd_data[31]) );
  OA21X1 U414 ( .A0(f32_mux_0_data[12]), .A1(f32_mux_1_data[12]), .B0(n337), .Y(o_rd_data[12]) );
  OA21X1 U415 ( .A0(f32_mux_0_data[17]), .A1(f32_mux_1_data[17]), .B0(n336), .Y(o_rd_data[17]) );
  OA21X1 U416 ( .A0(f32_mux_0_data[9]), .A1(f32_mux_1_data[9]), .B0(n336), .Y(o_rd_data[9]) );
  OA21X1 U417 ( .A0(f32_mux_0_data[10]), .A1(f32_mux_1_data[10]), .B0(n337), .Y(o_rd_data[10]) );
  OA21X1 U418 ( .A0(f32_mux_0_data[6]), .A1(f32_mux_1_data[6]), .B0(n337), .Y(o_rd_data[6]) );
  OA21X1 U419 ( .A0(f32_mux_0_data[15]), .A1(f32_mux_1_data[15]), .B0(n337), .Y(o_rd_data[15]) );
  OA21X1 U420 ( .A0(f32_mux_0_data[11]), .A1(f32_mux_1_data[11]), .B0(n336), .Y(o_rd_data[11]) );
  OA21X1 U421 ( .A0(f32_mux_0_data[1]), .A1(f32_mux_1_data[1]), .B0(n337), .Y(o_rd_data[1]) );
  OA21X1 U422 ( .A0(f32_mux_0_data[5]), .A1(f32_mux_1_data[5]), .B0(n337), .Y(o_rd_data[5]) );
  OA21X1 U423 ( .A0(f32_mux_0_data[8]), .A1(f32_mux_1_data[8]), .B0(n336), .Y(o_rd_data[8]) );
  OA21X1 U424 ( .A0(f32_mux_0_data[7]), .A1(f32_mux_1_data[7]), .B0(n337), .Y(o_rd_data[7]) );
  OA21X1 U425 ( .A0(f32_mux_0_data[13]), .A1(f32_mux_1_data[13]), .B0(n337), .Y(o_rd_data[13]) );
  AOI22X1 U426 ( .A0(n170), .A1(i_hisbuf0_3[17]), .B0(n168), .B1(i_hisbuf0_2[17]), .Y(n348) );
  AOI22X1 U427 ( .A0(n857), .A1(i_hisbuf2_2[17]), .B0(i_hisbuf1_2[17]), .B1(n166), .Y(n347) );
  AOI22X1 U428 ( .A0(n838), .A1(i_hisbuf1_0[17]), .B0(i_hisbuf2_0[17]), .B1(n830), .Y(n341) );
  AOI22X1 U429 ( .A0(n311), .A1(i_hisbuf0_1[17]), .B0(n816), .B1(i_hisbuf1_1[17]), .Y(n339) );
  AOI22X1 U430 ( .A0(n843), .A1(i_hisbuf3_1[17]), .B0(n130), .B1(i_spare_config[17]), .Y(n338) );
  NAND4X1 U431 ( .A(n341), .B(n340), .C(n339), .D(n338), .Y(n345) );
  INVX2 U432 ( .A(n159), .Y(n396) );
  AOI22X1 U433 ( .A0(n165), .A1(i_hisbuf1_3[17]), .B0(n821), .B1(i_hisbuf3_2[17]), .Y(n343) );
  AO21X1 U434 ( .A0(n823), .A1(i_hisbuf0_0[17]), .B0(n343_inv), .Y(n344) );
  AOI21X1 U435 ( .A0(n852), .A1(n345), .B0(n344), .Y(n346) );
  AOI22X1 U436 ( .A0(n170), .A1(i_hisbuf0_3[21]), .B0(n168), .B1(i_hisbuf0_2[21]), .Y(n358) );
  AOI22X1 U437 ( .A0(n857), .A1(i_hisbuf2_2[21]), .B0(i_hisbuf1_2[21]), .B1(n166), .Y(n357) );
  AOI22X1 U438 ( .A0(n838), .A1(i_hisbuf1_0[21]), .B0(i_hisbuf2_0[21]), .B1(n830), .Y(n352) );
  AOI22X1 U439 ( .A0(n815), .A1(i_hisbuf3_0[21]), .B0(n836), .B1(i_hisbuf2_1[21]), .Y(n351) );
  AOI22X1 U440 ( .A0(n311), .A1(i_hisbuf0_1[21]), .B0(n816), .B1(i_hisbuf1_1[21]), .Y(n350) );
  AOI22X1 U441 ( .A0(n843), .A1(i_hisbuf3_1[21]), .B0(n130), .B1(i_spare_config[21]), .Y(n349) );
  NAND4X1 U442 ( .A(n352), .B(n351), .C(n350), .D(n349), .Y(n355) );
  AOI22X1 U443 ( .A0(n165), .A1(i_hisbuf1_3[21]), .B0(n807), .B1(i_hisbuf3_2[21]), .Y(n353) );
  AOI21X1 U444 ( .A0(n852), .A1(n355), .B0(n354), .Y(n356) );
  AOI22X1 U445 ( .A0(n170), .A1(i_hisbuf0_3[22]), .B0(n168), .B1(i_hisbuf0_2[22]), .Y(n368) );
  AOI22X1 U446 ( .A0(n857), .A1(i_hisbuf2_2[22]), .B0(i_hisbuf1_2[22]), .B1(n166), .Y(n367) );
  AOI22X1 U447 ( .A0(n838), .A1(i_hisbuf1_0[22]), .B0(i_hisbuf2_0[22]), .B1(n830), .Y(n362) );
  AOI22X1 U448 ( .A0(n815), .A1(i_hisbuf3_0[22]), .B0(n836), .B1(i_hisbuf2_1[22]), .Y(n361) );
  AOI22X1 U449 ( .A0(n311), .A1(i_hisbuf0_1[22]), .B0(n816), .B1(i_hisbuf1_1[22]), .Y(n360) );
  AOI22X1 U450 ( .A0(n843), .A1(i_hisbuf3_1[22]), .B0(n130), .B1(i_spare_config[22]), .Y(n359) );
  NAND4X1 U451 ( .A(n362), .B(n361), .C(n360), .D(n359), .Y(n365) );
  AOI22X1 U452 ( .A0(n165), .A1(i_hisbuf1_3[22]), .B0(n807), .B1(i_hisbuf3_2[22]), .Y(n363) );
  AO21X1 U453 ( .A0(n823), .A1(i_hisbuf0_0[22]), .B0(n363_inv), .Y(n364) );
  AOI21X1 U454 ( .A0(n852), .A1(n365), .B0(n364), .Y(n366) );
  INVX2 U455 ( .A(n500), .Y(n597) );
  NAND3X2 U456 ( .A(n371), .B(n372), .C(scan_iso_or2), .Y(n394) );
  NOR2X4 U457 ( .A(n382), .B(n394), .Y(n657) );
  BUFX4 U458 ( .A(n736), .Y(n751) );
  AOI22X1 U459 ( .A0(n657), .A1(i_hisbuf1_4[23]), .B0(n751), .B1(i_hisbuf2_5[23]), .Y(n378) );
  NOR2X4 U460 ( .A(n380), .B(n394), .Y(n640) );
  NOR2X2 U461 ( .A(n386), .B(n394), .Y(n704) );
  NOR2X2 U462 ( .A(n386), .B(n373), .Y(n658) );
  BUFX4 U463 ( .A(n658), .Y(n753) );
  AOI22X1 U464 ( .A0(n753), .A1(i_hisbuf3_5[23]), .B0(n641), .B1(i_hisbuf0_6[23]), .Y(n376) );
  NOR2X4 U465 ( .A(n382), .B(n373), .Y(n642) );
  AND2X2 U466 ( .A(scan_iso_or5), .B(n374), .Y(n705) );
  AOI22X1 U467 ( .A0(n642), .A1(i_hisbuf1_6[23]), .B0(n705), .B1(i_hisbuf3_6[23]), .Y(n375) );
  NAND4X1 U468 ( .A(n378), .B(n377), .C(n376), .D(n375), .Y(n392) );
  NOR2X4 U469 ( .A(n380), .B(n381), .Y(n663) );
  AOI22X1 U470 ( .A0(n663), .A1(i_hisbuf0_5[23]), .B0(n710), .B1(i_hisbuf3_4[23]), .Y(n390) );
  NOR2X4 U471 ( .A(n382), .B(n381), .Y(n664) );
  AOI22X1 U472 ( .A0(n564), .A1(i_hisbuf0_7[23]), .B0(n664), .B1(i_hisbuf1_5[23]), .Y(n389) );
  NOR3X2 U473 ( .A(n395), .B(n383), .C(n393), .Y(n492) );
  AND2X2 U474 ( .B(n839), .A(n395_inv), .Y(n665) );
  INVX1 U474_inv ( .A(n395), .Y(n395_inv) );
  AOI22X1 U475 ( .A0(n666), .A1(i_hisbuf2_6[23]), .B0(n665), .B1(i_hisbuf2_7[23]), .Y(n388) );
  NOR2X4 U476 ( .A(n384), .B(n395), .Y(n667) );
  NOR3X2 U477 ( .A(n395), .B(n386), .C(n385), .Y(n711) );
  AOI22X1 U478 ( .A0(n667), .A1(i_hisbuf1_7[23]), .B0(n711), .B1(i_hisbuf3_7[23]), .Y(n387) );
  NAND4X1 U479 ( .A(n390), .B(n389), .C(n388), .D(n387), .Y(n391) );
  AOI21X1 U480 ( .A0(n597), .A1(n392), .B0(n391), .Y(n398) );
  NOR2X4 U481 ( .A(n396), .B(n395), .Y(n768) );
  BUFX6 U482 ( .A(n768), .Y(n732) );
  AOI22X1 U483 ( .A0(n674), .A1(i_hisbuf2_3[23]), .B0(n732), .B1(i_agg_su_count_a[23]), .Y(n397) );
  AOI22X1 U484 ( .A0(n657), .A1(i_hisbuf1_4[22]), .B0(n751), .B1(i_hisbuf2_5[22]), .Y(n403) );
  AOI22X1 U485 ( .A0(n640), .A1(i_hisbuf0_4[22]), .B0(n704), .B1(i_hisbuf3_3[22]), .Y(n402) );
  AOI22X1 U486 ( .A0(n658), .A1(i_hisbuf3_5[22]), .B0(n641), .B1(i_hisbuf0_6[22]), .Y(n401) );
  AOI22X1 U487 ( .A0(n642), .A1(i_hisbuf1_6[22]), .B0(n705), .B1(i_hisbuf3_6[22]), .Y(n400) );
  NAND4X1 U488 ( .A(n403), .B(n402), .C(n401), .D(n400), .Y(n409) );
  BUFX4 U489 ( .A(n710), .Y(n759) );
  AOI22X1 U490 ( .A0(n663), .A1(i_hisbuf0_5[22]), .B0(n759), .B1(i_hisbuf3_4[22]), .Y(n407) );
  AOI22X1 U491 ( .A0(n564), .A1(i_hisbuf0_7[22]), .B0(n664), .B1(i_hisbuf1_5[22]), .Y(n406) );
  AOI22X1 U492 ( .A0(n666), .A1(i_hisbuf2_6[22]), .B0(n665), .B1(i_hisbuf2_7[22]), .Y(n405) );
  AOI22X1 U493 ( .A0(n667), .A1(i_hisbuf1_7[22]), .B0(n711), .B1(i_hisbuf3_7[22]), .Y(n404) );
  NAND4X1 U494 ( .A(n407), .B(n406), .C(n405), .D(n404), .Y(n408) );
  AOI21X1 U495 ( .A0(n597), .A1(n409), .B0(n408), .Y(n411) );
  AOI22X1 U496 ( .A0(n674), .A1(i_hisbuf2_3[22]), .B0(n732), .B1(i_agg_su_count_a[22]), .Y(n410) );
  AOI22X1 U497 ( .A0(n657), .A1(i_hisbuf1_4[6]), .B0(n751), .B1(i_hisbuf2_5[6]), .Y(n416) );
  AOI22X1 U498 ( .A0(n640), .A1(i_hisbuf0_4[6]), .B0(n704), .B1(i_hisbuf3_3[6]), .Y(n415) );
  AOI22X1 U499 ( .A0(n658), .A1(i_hisbuf3_5[6]), .B0(n641), .B1(i_hisbuf0_6[6]), .Y(n414) );
  NAND4X1 U500 ( .A(n416), .B(n415), .C(n414), .D(n413), .Y(n422) );
  AOI22X1 U501 ( .A0(n663), .A1(i_hisbuf0_5[6]), .B0(n759), .B1(i_hisbuf3_4[6]), .Y(n420) );
  AOI22X1 U502 ( .A0(n564), .A1(i_hisbuf0_7[6]), .B0(n664), .B1(i_hisbuf1_5[6]), .Y(n419) );
  AOI22X1 U503 ( .A0(n666), .A1(i_hisbuf2_6[6]), .B0(n665), .B1(i_hisbuf2_7[6]), .Y(n418) );
  AOI22X1 U504 ( .A0(n667), .A1(i_hisbuf1_7[6]), .B0(n711), .B1(i_hisbuf3_7[6]), .Y(n417) );
  NAND4X1 U505 ( .A(n420), .B(n419), .C(n418), .D(n417), .Y(n421) );
  AOI21X1 U506 ( .A0(n597), .A1(n422), .B0(n421), .Y(n424) );
  AOI22X1 U507 ( .A0(n674), .A1(i_hisbuf2_3[6]), .B0(n732), .B1(i_agg_su_count_a[6]), .Y(n423) );
  AOI22X1 U508 ( .A0(n657), .A1(i_hisbuf1_4[7]), .B0(n751), .B1(i_hisbuf2_5[7]), .Y(n429) );
  AOI22X1 U509 ( .A0(n640), .A1(i_hisbuf0_4[7]), .B0(n704), .B1(i_hisbuf3_3[7]), .Y(n428) );
  AOI22X1 U510 ( .A0(n658), .A1(i_hisbuf3_5[7]), .B0(n641), .B1(i_hisbuf0_6[7]), .Y(n427) );
  AOI22X1 U511 ( .A0(n642), .A1(i_hisbuf1_6[7]), .B0(n705), .B1(i_hisbuf3_6[7]), .Y(n426) );
  NAND4X1 U512 ( .A(n429), .B(n428), .C(n427), .D(n426), .Y(n435) );
  AOI22X1 U513 ( .A0(n663), .A1(i_hisbuf0_5[7]), .B0(n759), .B1(i_hisbuf3_4[7]), .Y(n433) );
  AOI22X1 U514 ( .A0(n564), .A1(i_hisbuf0_7[7]), .B0(n664), .B1(i_hisbuf1_5[7]), .Y(n432) );
  AOI22X1 U515 ( .A0(n666), .A1(i_hisbuf2_6[7]), .B0(n665), .B1(i_hisbuf2_7[7]), .Y(n431) );
  AOI22X1 U516 ( .A0(n667), .A1(i_hisbuf1_7[7]), .B0(n711), .B1(i_hisbuf3_7[7]), .Y(n430) );
  NAND4X1 U517 ( .A(n433), .B(n432), .C(n431), .D(n430), .Y(n434) );
  AOI21X1 U518 ( .A0(n597), .A1(n435), .B0(n434), .Y(n437) );
  AOI22X1 U519 ( .A0(n674), .A1(i_hisbuf2_3[7]), .B0(n732), .B1(i_agg_su_count_a[7]), .Y(n436) );
  NAND2X1 U520 ( .A(n656), .B(i_hisbuf2_4[1]), .Y(n451) );
  AOI22X1 U521 ( .A0(n657), .A1(i_hisbuf1_4[1]), .B0(n751), .B1(i_hisbuf2_5[1]), .Y(n442) );
  AOI22X1 U522 ( .A0(n658), .A1(i_hisbuf3_5[1]), .B0(n641), .B1(i_hisbuf0_6[1]), .Y(n440) );
  AOI22X1 U523 ( .A0(n642), .A1(i_hisbuf1_6[1]), .B0(n705), .B1(i_hisbuf3_6[1]), .Y(n439) );
  NAND4X1 U524 ( .A(n442), .B(n441), .C(n440), .D(n439), .Y(n448) );
  AOI22X1 U525 ( .A0(n663), .A1(i_hisbuf0_5[1]), .B0(n759), .B1(i_hisbuf3_4[1]), .Y(n446) );
  AOI22X1 U526 ( .A0(n564), .A1(i_hisbuf0_7[1]), .B0(n664), .B1(i_hisbuf1_5[1]), .Y(n445) );
  AOI22X1 U527 ( .A0(n666), .A1(i_hisbuf2_6[1]), .B0(n665), .B1(i_hisbuf2_7[1]), .Y(n444) );
  AOI22X1 U528 ( .A0(n667), .A1(i_hisbuf1_7[1]), .B0(n711), .B1(i_hisbuf3_7[1]), .Y(n443) );
  NAND4X1 U529 ( .A(n446), .B(n445), .C(n444), .D(n443), .Y(n447) );
  AOI21X1 U530 ( .A0(n597), .A1(n448), .B0(n447), .Y(n450) );
  AOI22X1 U531 ( .A0(n769), .A1(i_hisbuf2_3[1]), .B0(n768), .B1(i_agg_su_count_a[1]), .Y(n449) );
  AOI22X1 U532 ( .A0(n656), .A1(i_hisbuf2_4[30]), .B0(n769), .B1(i_hisbuf2_3[30]), .Y(n454) );
  AND2X1 U533 ( .B(n751), .A(n500_inv), .Y(n474) );
  INVX1 U533_inv ( .A(n500), .Y(n500_inv) );
  AOI22X1 U534 ( .A0(n492), .A1(i_hisbuf2_6[30]), .B0(i_hisbuf2_5[30]), .B1(n474), .Y(n453) );
  AOI22X1 U535 ( .A0(n768), .A1(i_agg_su_count_a[30]), .B0(n665), .B1(i_hisbuf2_7[30]), .Y(n452) );
  AOI22X1 U536 ( .A0(n657), .A1(i_hisbuf1_4[8]), .B0(n751), .B1(i_hisbuf2_5[8]), .Y(n458) );
  BUFX4 U537 ( .A(n704), .Y(n752) );
  AOI22X1 U538 ( .A0(n753), .A1(i_hisbuf3_5[8]), .B0(n641), .B1(i_hisbuf0_6[8]), .Y(n456) );
  AOI22X1 U539 ( .A0(n642), .A1(i_hisbuf1_6[8]), .B0(n705), .B1(i_hisbuf3_6[8]), .Y(n455) );
  NAND4X1 U540 ( .A(n458), .B(n457), .C(n456), .D(n455), .Y(n464) );
  AOI22X1 U541 ( .A0(n663), .A1(i_hisbuf0_5[8]), .B0(n759), .B1(i_hisbuf3_4[8]), .Y(n462) );
  AOI22X1 U542 ( .A0(n564), .A1(i_hisbuf0_7[8]), .B0(n664), .B1(i_hisbuf1_5[8]), .Y(n461) );
  AOI22X1 U543 ( .A0(n666), .A1(i_hisbuf2_6[8]), .B0(n665), .B1(i_hisbuf2_7[8]), .Y(n460) );
  AOI22X1 U544 ( .A0(n667), .A1(i_hisbuf1_7[8]), .B0(n711), .B1(i_hisbuf3_7[8]), .Y(n459) );
  NAND4X1 U545 ( .A(n462), .B(n461), .C(n460), .D(n459), .Y(n463) );
  AOI21X1 U546 ( .A0(n597), .A1(n464), .B0(n463), .Y(n466) );
  AOI22X1 U547 ( .A0(n769), .A1(i_hisbuf2_3[8]), .B0(n768), .B1(i_agg_su_count_a[8]), .Y(n465) );
  AOI22X1 U548 ( .A0(n656), .A1(i_hisbuf2_4[28]), .B0(n674), .B1(i_hisbuf2_3[28]), .Y(n470) );
  AOI22X1 U549 ( .A0(n666), .A1(i_hisbuf2_6[28]), .B0(i_hisbuf2_5[28]), .B1(n474), .Y(n469) );
  BUFX4 U550 ( .A(n665), .Y(n760) );
  AOI22X1 U551 ( .A0(n732), .A1(i_agg_su_count_a[28]), .B0(n760), .B1(i_hisbuf2_7[28]), .Y(n468) );
  AOI22X1 U552 ( .A0(n656), .A1(i_hisbuf2_4[29]), .B0(n674), .B1(i_hisbuf2_3[29]), .Y(n473) );
  AOI22X1 U553 ( .A0(n492), .A1(i_hisbuf2_6[29]), .B0(i_hisbuf2_5[29]), .B1(n474), .Y(n472) );
  AOI22X1 U554 ( .A0(n656), .A1(i_hisbuf2_4[27]), .B0(n674), .B1(i_hisbuf2_3[27]), .Y(n477) );
  AOI22X1 U555 ( .A0(n492), .A1(i_hisbuf2_6[27]), .B0(i_hisbuf2_5[27]), .B1(n474), .Y(n476) );
  AOI22X1 U556 ( .A0(n768), .A1(i_agg_su_count_a[27]), .B0(n665), .B1(i_hisbuf2_7[27]), .Y(n475) );
  AOI22X1 U557 ( .A0(n710), .A1(i_hisbuf3_4[25]), .B0(i_hisbuf3_7[25]), .B1(n761), .Y(n484) );
  AOI22X1 U558 ( .A0(n492), .A1(i_hisbuf2_6[25]), .B0(n665), .B1(i_hisbuf2_7[25]), .Y(n483) );
  AOI22X1 U559 ( .A0(n751), .A1(i_hisbuf2_5[25]), .B0(i_hisbuf3_3[25]), .B1(n752), .Y(n479) );
  AOI22X1 U560 ( .A0(n753), .A1(i_hisbuf3_5[25]), .B0(i_hisbuf3_6[25]), .B1(n705), .Y(n478) );
  AOI21X1 U561 ( .A0(n479), .A1(n478), .B0(n500), .Y(n480) );
  AOI211X1 U562 ( .A0(i_hisbuf2_4[25]), .A1(n656), .B0(n481), .C0(n480), .Y(n482) );
  AOI22X1 U563 ( .A0(n710), .A1(i_hisbuf3_4[26]), .B0(i_hisbuf3_7[26]), .B1(n761), .Y(n491) );
  AOI22X1 U564 ( .A0(n492), .A1(i_hisbuf2_6[26]), .B0(n665), .B1(i_hisbuf2_7[26]), .Y(n490) );
  AOI22X1 U565 ( .A0(n753), .A1(i_hisbuf3_5[26]), .B0(i_hisbuf3_6[26]), .B1(n705), .Y(n485) );
  AOI21X1 U566 ( .A0(n486), .A1(n485), .B0(n500), .Y(n487) );
  AOI211X1 U567 ( .A0(i_hisbuf2_4[26]), .A1(n656), .B0(n488), .C0(n487), .Y(n489) );
  AOI22X1 U568 ( .A0(n710), .A1(i_hisbuf3_4[24]), .B0(i_hisbuf3_7[24]), .B1(n761), .Y(n499) );
  AOI22X1 U569 ( .A0(n492), .A1(i_hisbuf2_6[24]), .B0(n665), .B1(i_hisbuf2_7[24]), .Y(n498) );
  AOI22X1 U570 ( .A0(n751), .A1(i_hisbuf2_5[24]), .B0(i_hisbuf3_3[24]), .B1(n752), .Y(n494) );
  AOI22X1 U571 ( .A0(n658), .A1(i_hisbuf3_5[24]), .B0(i_hisbuf3_6[24]), .B1(n705), .Y(n493) );
  AOI21X1 U572 ( .A0(n494), .A1(n493), .B0(n500), .Y(n495) );
  AOI211X1 U573 ( .A0(i_hisbuf2_4[24]), .A1(n656), .B0(n496), .C0(n495), .Y(n497) );
  AOI22X1 U574 ( .A0(n710), .A1(i_hisbuf3_4[27]), .B0(i_hisbuf3_7[27]), .B1(n761), .Y(n507) );
  AOI22X1 U575 ( .A0(n666), .A1(i_hisbuf2_6[31]), .B0(n665), .B1(i_hisbuf2_7[31]), .Y(n506) );
  AOI22X1 U576 ( .A0(n751), .A1(i_hisbuf2_5[31]), .B0(i_hisbuf3_3[27]), .B1(n704), .Y(n502) );
  AOI22X1 U577 ( .A0(n753), .A1(i_hisbuf3_5[27]), .B0(i_hisbuf3_6[27]), .B1(n705), .Y(n501) );
  AOI21X1 U578 ( .A0(n502), .A1(n501), .B0(n500), .Y(n503) );
  AOI211X1 U579 ( .A0(i_hisbuf2_4[31]), .A1(n656), .B0(n504), .C0(n503), .Y(n505) );
  AOI22X1 U580 ( .A0(n657), .A1(i_hisbuf1_4[19]), .B0(n751), .B1(i_hisbuf2_5[19]), .Y(n511) );
  AOI22X1 U581 ( .A0(n640), .A1(i_hisbuf0_4[19]), .B0(n752), .B1(i_hisbuf3_3[19]), .Y(n510) );
  AOI22X1 U582 ( .A0(n753), .A1(i_hisbuf3_5[19]), .B0(n641), .B1(i_hisbuf0_6[19]), .Y(n509) );
  NAND4X1 U583 ( .A(n511), .B(n510), .C(n509), .D(n508), .Y(n517) );
  AOI22X1 U584 ( .A0(n663), .A1(i_hisbuf0_5[19]), .B0(n759), .B1(i_hisbuf3_4[19]), .Y(n515) );
  AOI22X1 U585 ( .A0(n564), .A1(i_hisbuf0_7[19]), .B0(n664), .B1(i_hisbuf1_5[19]), .Y(n514) );
  AOI22X1 U586 ( .A0(n492), .A1(i_hisbuf2_6[19]), .B0(n665), .B1(i_hisbuf2_7[19]), .Y(n513) );
  AOI22X1 U587 ( .A0(n667), .A1(i_hisbuf1_7[19]), .B0(n761), .B1(i_hisbuf3_7[19]), .Y(n512) );
  NAND4X1 U588 ( .A(n515), .B(n514), .C(n513), .D(n512), .Y(n516) );
  AOI21X1 U589 ( .A0(n597), .A1(n517), .B0(n516), .Y(n519) );
  AOI22X1 U590 ( .A0(n657), .A1(i_hisbuf1_4[18]), .B0(n736), .B1(i_hisbuf2_5[18]), .Y(n524) );
  AOI22X1 U591 ( .A0(n640), .A1(i_hisbuf0_4[18]), .B0(n752), .B1(i_hisbuf3_3[18]), .Y(n523) );
  AOI22X1 U592 ( .A0(n753), .A1(i_hisbuf3_5[18]), .B0(n641), .B1(i_hisbuf0_6[18]), .Y(n522) );
  BUFX4 U593 ( .A(n705), .Y(n754) );
  AOI22X1 U594 ( .A0(n642), .A1(i_hisbuf1_6[18]), .B0(n754), .B1(i_hisbuf3_6[18]), .Y(n521) );
  NAND4X1 U595 ( .A(n524), .B(n523), .C(n522), .D(n521), .Y(n530) );
  AOI22X1 U596 ( .A0(n663), .A1(i_hisbuf0_5[18]), .B0(n759), .B1(i_hisbuf3_4[18]), .Y(n528) );
  AOI22X1 U597 ( .A0(n564), .A1(i_hisbuf0_7[18]), .B0(n664), .B1(i_hisbuf1_5[18]), .Y(n527) );
  AOI22X1 U598 ( .A0(n666), .A1(i_hisbuf2_6[18]), .B0(n665), .B1(i_hisbuf2_7[18]), .Y(n526) );
  AOI22X1 U599 ( .A0(n667), .A1(i_hisbuf1_7[18]), .B0(n761), .B1(i_hisbuf3_7[18]), .Y(n525) );
  NAND4X1 U600 ( .A(n528), .B(n527), .C(n526), .D(n525), .Y(n529) );
  AOI21X1 U601 ( .A0(n597), .A1(n530), .B0(n529), .Y(n532) );
  AOI22X1 U602 ( .A0(n769), .A1(i_hisbuf2_3[18]), .B0(n768), .B1(i_agg_su_count_a[18]), .Y(n531) );
  AOI22X1 U603 ( .A0(n657), .A1(i_hisbuf1_4[20]), .B0(n751), .B1(i_hisbuf2_5[20]), .Y(n537) );
  AOI22X1 U604 ( .A0(n640), .A1(i_hisbuf0_4[20]), .B0(n704), .B1(i_hisbuf3_3[20]), .Y(n536) );
  AOI22X1 U605 ( .A0(n753), .A1(i_hisbuf3_5[20]), .B0(n641), .B1(i_hisbuf0_6[20]), .Y(n535) );
  AOI22X1 U606 ( .A0(n642), .A1(i_hisbuf1_6[20]), .B0(n754), .B1(i_hisbuf3_6[20]), .Y(n534) );
  NAND4X1 U607 ( .A(n537), .B(n536), .C(n535), .D(n534), .Y(n543) );
  AOI22X1 U608 ( .A0(n663), .A1(i_hisbuf0_5[20]), .B0(n759), .B1(i_hisbuf3_4[20]), .Y(n541) );
  AOI22X1 U609 ( .A0(n564), .A1(i_hisbuf0_7[20]), .B0(n664), .B1(i_hisbuf1_5[20]), .Y(n540) );
  AOI22X1 U610 ( .A0(n666), .A1(i_hisbuf2_6[20]), .B0(n665), .B1(i_hisbuf2_7[20]), .Y(n539) );
  AOI22X1 U611 ( .A0(n667), .A1(i_hisbuf1_7[20]), .B0(n761), .B1(i_hisbuf3_7[20]), .Y(n538) );
  NAND4X1 U612 ( .A(n541), .B(n540), .C(n539), .D(n538), .Y(n542) );
  AOI21X1 U613 ( .A0(n597), .A1(n543), .B0(n542), .Y(n545) );
  AOI22X1 U614 ( .A0(n674), .A1(i_hisbuf2_3[20]), .B0(n732), .B1(i_agg_su_count_a[20]), .Y(n544) );
  AOI22X1 U615 ( .A0(n657), .A1(i_hisbuf1_4[21]), .B0(n751), .B1(i_hisbuf2_5[21]), .Y(n550) );
  AOI22X1 U616 ( .A0(n640), .A1(i_hisbuf0_4[21]), .B0(n704), .B1(i_hisbuf3_3[21]), .Y(n549) );
  AOI22X1 U617 ( .A0(n642), .A1(i_hisbuf1_6[21]), .B0(n705), .B1(i_hisbuf3_6[21]), .Y(n547) );
  NAND4X1 U618 ( .A(n550), .B(n549), .C(n548), .D(n547), .Y(n556) );
  AOI22X1 U619 ( .A0(n663), .A1(i_hisbuf0_5[21]), .B0(n759), .B1(i_hisbuf3_4[21]), .Y(n554) );
  AOI22X1 U620 ( .A0(n564), .A1(i_hisbuf0_7[21]), .B0(n664), .B1(i_hisbuf1_5[21]), .Y(n553) );
  AOI22X1 U621 ( .A0(n666), .A1(i_hisbuf2_6[21]), .B0(n665), .B1(i_hisbuf2_7[21]), .Y(n552) );
  AOI22X1 U622 ( .A0(n667), .A1(i_hisbuf1_7[21]), .B0(n761), .B1(i_hisbuf3_7[21]), .Y(n551) );
  NAND4X1 U623 ( .A(n554), .B(n553), .C(n552), .D(n551), .Y(n555) );
  AOI21X1 U624 ( .A0(n597), .A1(n556), .B0(n555), .Y(n558) );
  AOI22X1 U625 ( .A0(n674), .A1(i_hisbuf2_3[21]), .B0(n732), .B1(i_agg_su_count_a[21]), .Y(n557) );
  AOI22X1 U626 ( .A0(n657), .A1(i_hisbuf1_4[17]), .B0(n736), .B1(i_hisbuf2_5[17]), .Y(n563) );
  AOI22X1 U627 ( .A0(n640), .A1(i_hisbuf0_4[17]), .B0(n752), .B1(i_hisbuf3_3[17]), .Y(n562) );
  AOI22X1 U628 ( .A0(n753), .A1(i_hisbuf3_5[17]), .B0(n641), .B1(i_hisbuf0_6[17]), .Y(n561) );
  AOI22X1 U629 ( .A0(n642), .A1(i_hisbuf1_6[17]), .B0(n754), .B1(i_hisbuf3_6[17]), .Y(n560) );
  NAND4X1 U630 ( .A(n563), .B(n562), .C(n561), .D(n560), .Y(n570) );
  AOI22X1 U631 ( .A0(n564), .A1(i_hisbuf0_7[17]), .B0(n664), .B1(i_hisbuf1_5[17]), .Y(n567) );
  AOI22X1 U632 ( .A0(n666), .A1(i_hisbuf2_6[17]), .B0(n760), .B1(i_hisbuf2_7[17]), .Y(n566) );
  AOI22X1 U633 ( .A0(n667), .A1(i_hisbuf1_7[17]), .B0(n761), .B1(i_hisbuf3_7[17]), .Y(n565) );
  NAND4X1 U634 ( .A(n568), .B(n567), .C(n566), .D(n565), .Y(n569) );
  AOI21X1 U635 ( .A0(n597), .A1(n570), .B0(n569), .Y(n572) );
  AOI22X1 U636 ( .A0(n769), .A1(i_hisbuf2_3[17]), .B0(n768), .B1(i_agg_su_count_a[17]), .Y(n571) );
  AOI22X1 U637 ( .A0(n657), .A1(i_hisbuf1_4[16]), .B0(n736), .B1(i_hisbuf2_5[16]), .Y(n577) );
  AOI22X1 U638 ( .A0(n640), .A1(i_hisbuf0_4[16]), .B0(n752), .B1(i_hisbuf3_3[16]), .Y(n576) );
  AOI22X1 U639 ( .A0(n753), .A1(i_hisbuf3_5[16]), .B0(n641), .B1(i_hisbuf0_6[16]), .Y(n575) );
  AOI22X1 U640 ( .A0(n642), .A1(i_hisbuf1_6[16]), .B0(n754), .B1(i_hisbuf3_6[16]), .Y(n574) );
  NAND4X1 U641 ( .A(n577), .B(n576), .C(n575), .D(n574), .Y(n583) );
  AOI22X1 U642 ( .A0(n663), .A1(i_hisbuf0_5[16]), .B0(n759), .B1(i_hisbuf3_4[16]), .Y(n581) );
  AOI22X1 U643 ( .A0(n564), .A1(i_hisbuf0_7[16]), .B0(n664), .B1(i_hisbuf1_5[16]), .Y(n580) );
  AOI22X1 U644 ( .A0(n492), .A1(i_hisbuf2_6[16]), .B0(n760), .B1(i_hisbuf2_7[16]), .Y(n579) );
  AOI22X1 U645 ( .A0(n667), .A1(i_hisbuf1_7[16]), .B0(n761), .B1(i_hisbuf3_7[16]), .Y(n578) );
  NAND4X1 U646 ( .A(n581), .B(n580), .C(n579), .D(n578), .Y(n582) );
  AOI21X1 U647 ( .A0(n597), .A1(n583), .B0(n582), .Y(n585) );
  AOI22X1 U648 ( .A0(n769), .A1(i_hisbuf2_3[16]), .B0(n768), .B1(i_agg_su_count_a[16]), .Y(n584) );
  AOI22X1 U649 ( .A0(n657), .A1(i_hisbuf1_4[15]), .B0(n736), .B1(i_hisbuf2_5[15]), .Y(n590) );
  AOI22X1 U650 ( .A0(n640), .A1(i_hisbuf0_4[15]), .B0(n752), .B1(i_hisbuf3_3[15]), .Y(n589) );
  AOI22X1 U651 ( .A0(n753), .A1(i_hisbuf3_5[15]), .B0(n641), .B1(i_hisbuf0_6[15]), .Y(n588) );
  AOI22X1 U652 ( .A0(n642), .A1(i_hisbuf1_6[15]), .B0(n754), .B1(i_hisbuf3_6[15]), .Y(n587) );
  NAND4X1 U653 ( .A(n590), .B(n589), .C(n588), .D(n587), .Y(n596) );
  AOI22X1 U654 ( .A0(n663), .A1(i_hisbuf0_5[15]), .B0(n759), .B1(i_hisbuf3_4[15]), .Y(n594) );
  AOI22X1 U655 ( .A0(n666), .A1(i_hisbuf2_6[15]), .B0(n760), .B1(i_hisbuf2_7[15]), .Y(n592) );
  AOI22X1 U656 ( .A0(n667), .A1(i_hisbuf1_7[15]), .B0(n761), .B1(i_hisbuf3_7[15]), .Y(n591) );
  NAND4X1 U657 ( .A(n594), .B(n593), .C(n592), .D(n591), .Y(n595) );
  AOI21X1 U658 ( .A0(n597), .A1(n596), .B0(n595), .Y(n599) );
  AOI22X1 U659 ( .A0(n769), .A1(i_hisbuf2_3[15]), .B0(n732), .B1(i_agg_su_count_a[15]), .Y(n598) );
  AOI22X1 U660 ( .A0(n657), .A1(i_hisbuf1_4[0]), .B0(n736), .B1(i_hisbuf2_5[0]), .Y(n604) );
  AOI22X1 U661 ( .A0(n640), .A1(i_hisbuf0_4[0]), .B0(n752), .B1(i_hisbuf3_3[0]), .Y(n603) );
  AOI22X1 U662 ( .A0(n753), .A1(i_hisbuf3_5[0]), .B0(n641), .B1(i_hisbuf0_6[0]), .Y(n602) );
  AOI22X1 U663 ( .A0(n642), .A1(i_hisbuf1_6[0]), .B0(n705), .B1(i_hisbuf3_6[0]), .Y(n601) );
  NAND4X1 U664 ( .A(n604), .B(n603), .C(n602), .D(n601), .Y(n610) );
  AOI22X1 U665 ( .A0(n663), .A1(i_hisbuf0_5[0]), .B0(n710), .B1(i_hisbuf3_4[0]), .Y(n608) );
  AOI22X1 U666 ( .A0(n564), .A1(i_hisbuf0_7[0]), .B0(n664), .B1(i_hisbuf1_5[0]), .Y(n607) );
  AOI22X1 U667 ( .A0(n666), .A1(i_hisbuf2_6[0]), .B0(n665), .B1(i_hisbuf2_7[0]), .Y(n606) );
  AOI22X1 U668 ( .A0(n667), .A1(i_hisbuf1_7[0]), .B0(n761), .B1(i_hisbuf3_7[0]), .Y(n605) );
  NAND4X1 U669 ( .A(n608), .B(n607), .C(n606), .D(n605), .Y(n609) );
  AOI21X1 U670 ( .A0(n131), .A1(n610), .B0(n609), .Y(n612) );
  AOI22X1 U671 ( .A0(n769), .A1(i_hisbuf2_3[0]), .B0(n768), .B1(i_agg_su_count_a[0]), .Y(n611) );
  NAND2X1 U672 ( .A(n656), .B(i_hisbuf2_4[5]), .Y(n626) );
  AOI22X1 U673 ( .A0(n657), .A1(i_hisbuf1_4[5]), .B0(n751), .B1(i_hisbuf2_5[5]), .Y(n617) );
  AOI22X1 U674 ( .A0(n640), .A1(i_hisbuf0_4[5]), .B0(n752), .B1(i_hisbuf3_3[5]), .Y(n616) );
  AOI22X1 U675 ( .A0(n658), .A1(i_hisbuf3_5[5]), .B0(n641), .B1(i_hisbuf0_6[5]), .Y(n615) );
  AOI22X1 U676 ( .A0(n642), .A1(i_hisbuf1_6[5]), .B0(n705), .B1(i_hisbuf3_6[5]), .Y(n614) );
  NAND4X1 U677 ( .A(n617), .B(n616), .C(n615), .D(n614), .Y(n623) );
  AOI22X1 U678 ( .A0(n663), .A1(i_hisbuf0_5[5]), .B0(n759), .B1(i_hisbuf3_4[5]), .Y(n621) );
  AOI22X1 U679 ( .A0(n564), .A1(i_hisbuf0_7[5]), .B0(n664), .B1(i_hisbuf1_5[5]), .Y(n620) );
  AOI22X1 U680 ( .A0(n666), .A1(i_hisbuf2_6[5]), .B0(n665), .B1(i_hisbuf2_7[5]), .Y(n619) );
  AOI22X1 U681 ( .A0(n667), .A1(i_hisbuf1_7[5]), .B0(n761), .B1(i_hisbuf3_7[5]), .Y(n618) );
  NAND4X1 U682 ( .A(n621), .B(n620), .C(n619), .D(n618), .Y(n622) );
  AOI21X1 U683 ( .A0(n131), .A1(n623), .B0(n622), .Y(n625) );
  AOI22X1 U684 ( .A0(n769), .A1(i_hisbuf2_3[5]), .B0(n768), .B1(i_agg_su_count_a[5]), .Y(n624) );
  AOI22X1 U685 ( .A0(n657), .A1(i_hisbuf1_4[3]), .B0(n751), .B1(i_hisbuf2_5[3]), .Y(n630) );
  AOI22X1 U686 ( .A0(n640), .A1(i_hisbuf0_4[3]), .B0(n752), .B1(i_hisbuf3_3[3]), .Y(n629) );
  AOI22X1 U687 ( .A0(n658), .A1(i_hisbuf3_5[3]), .B0(n641), .B1(i_hisbuf0_6[3]), .Y(n628) );
  AOI22X1 U688 ( .A0(n642), .A1(i_hisbuf1_6[3]), .B0(n705), .B1(i_hisbuf3_6[3]), .Y(n627) );
  NAND4X1 U689 ( .A(n630), .B(n629), .C(n628), .D(n627), .Y(n636) );
  AOI22X1 U690 ( .A0(n663), .A1(i_hisbuf0_5[3]), .B0(n759), .B1(i_hisbuf3_4[3]), .Y(n634) );
  AOI22X1 U691 ( .A0(n564), .A1(i_hisbuf0_7[3]), .B0(n664), .B1(i_hisbuf1_5[3]), .Y(n633) );
  AOI22X1 U692 ( .A0(n666), .A1(i_hisbuf2_6[3]), .B0(n665), .B1(i_hisbuf2_7[3]), .Y(n632) );
  AOI22X1 U693 ( .A0(n667), .A1(i_hisbuf1_7[3]), .B0(n761), .B1(i_hisbuf3_7[3]), .Y(n631) );
  NAND4X1 U694 ( .A(n634), .B(n633), .C(n632), .D(n631), .Y(n635) );
  AOI21X1 U695 ( .A0(n131), .A1(n636), .B0(n635), .Y(n638) );
  AOI22X1 U696 ( .A0(n769), .A1(i_hisbuf2_3[3]), .B0(n768), .B1(i_agg_su_count_a[3]), .Y(n637) );
  AOI22X1 U697 ( .A0(n657), .A1(i_hisbuf1_4[2]), .B0(n751), .B1(i_hisbuf2_5[2]), .Y(n646) );
  AOI22X1 U698 ( .A0(n640), .A1(i_hisbuf0_4[2]), .B0(n752), .B1(i_hisbuf3_3[2]), .Y(n645) );
  AOI22X1 U699 ( .A0(n658), .A1(i_hisbuf3_5[2]), .B0(n641), .B1(i_hisbuf0_6[2]), .Y(n644) );
  AOI22X1 U700 ( .A0(n642), .A1(i_hisbuf1_6[2]), .B0(n705), .B1(i_hisbuf3_6[2]), .Y(n643) );
  NAND4X1 U701 ( .A(n646), .B(n645), .C(n644), .D(n643), .Y(n652) );
  AOI22X1 U702 ( .A0(n663), .A1(i_hisbuf0_5[2]), .B0(n759), .B1(i_hisbuf3_4[2]), .Y(n650) );
  AOI22X1 U703 ( .A0(n564), .A1(i_hisbuf0_7[2]), .B0(n664), .B1(i_hisbuf1_5[2]), .Y(n649) );
  AOI22X1 U704 ( .A0(n666), .A1(i_hisbuf2_6[2]), .B0(n665), .B1(i_hisbuf2_7[2]), .Y(n648) );
  AOI22X1 U705 ( .A0(n667), .A1(i_hisbuf1_7[2]), .B0(n761), .B1(i_hisbuf3_7[2]), .Y(n647) );
  NAND4X1 U706 ( .A(n650), .B(n649), .C(n648), .D(n647), .Y(n651) );
  AOI21X1 U707 ( .A0(n131), .A1(n652), .B0(n651), .Y(n654) );
  AOI22X1 U708 ( .A0(n769), .A1(i_hisbuf2_3[2]), .B0(n732), .B1(i_agg_su_count_a[2]), .Y(n653) );
  AOI22X1 U709 ( .A0(n657), .A1(i_hisbuf1_4[4]), .B0(n751), .B1(i_hisbuf2_5[4]), .Y(n662) );
  AOI22X1 U710 ( .A0(n640), .A1(i_hisbuf0_4[4]), .B0(n752), .B1(i_hisbuf3_3[4]), .Y(n661) );
  AOI22X1 U711 ( .A0(n658), .A1(i_hisbuf3_5[4]), .B0(n641), .B1(i_hisbuf0_6[4]), .Y(n660) );
  AOI22X1 U712 ( .A0(n642), .A1(i_hisbuf1_6[4]), .B0(n705), .B1(i_hisbuf3_6[4]), .Y(n659) );
  NAND4X1 U713 ( .A(n662), .B(n661), .C(n660), .D(n659), .Y(n673) );
  AOI22X1 U714 ( .A0(n663), .A1(i_hisbuf0_5[4]), .B0(n759), .B1(i_hisbuf3_4[4]), .Y(n671) );
  AOI22X1 U715 ( .A0(n666), .A1(i_hisbuf2_6[4]), .B0(n665), .B1(i_hisbuf2_7[4]), .Y(n669) );
  AOI22X1 U716 ( .A0(n667), .A1(i_hisbuf1_7[4]), .B0(n761), .B1(i_hisbuf3_7[4]), .Y(n668) );
  NAND4X1 U717 ( .A(n671), .B(n670), .C(n669), .D(n668), .Y(n672) );
  AOI21X1 U718 ( .A0(n597), .A1(n673), .B0(n672), .Y(n676) );
  AOI22X1 U719 ( .A0(n674), .A1(i_hisbuf2_3[4]), .B0(n732), .B1(i_agg_su_count_a[4]), .Y(n675) );
  AOI22X1 U720 ( .A0(n657), .A1(i_hisbuf1_4[14]), .B0(n736), .B1(i_hisbuf2_5[14]), .Y(n681) );
  AOI22X1 U721 ( .A0(n640), .A1(i_hisbuf0_4[14]), .B0(n752), .B1(i_hisbuf3_3[14]), .Y(n680) );
  AOI22X1 U722 ( .A0(n753), .A1(i_hisbuf3_5[14]), .B0(n641), .B1(i_hisbuf0_6[14]), .Y(n679) );
  AOI22X1 U723 ( .A0(n642), .A1(i_hisbuf1_6[14]), .B0(n754), .B1(i_hisbuf3_6[14]), .Y(n678) );
  NAND4X1 U724 ( .A(n681), .B(n680), .C(n679), .D(n678), .Y(n687) );
  AOI22X1 U725 ( .A0(n663), .A1(i_hisbuf0_5[14]), .B0(n759), .B1(i_hisbuf3_4[14]), .Y(n685) );
  AOI22X1 U726 ( .A0(n564), .A1(i_hisbuf0_7[14]), .B0(n664), .B1(i_hisbuf1_5[14]), .Y(n684) );
  AOI22X1 U727 ( .A0(n666), .A1(i_hisbuf2_6[14]), .B0(n760), .B1(i_hisbuf2_7[14]), .Y(n683) );
  AOI22X1 U728 ( .A0(n667), .A1(i_hisbuf1_7[14]), .B0(n761), .B1(i_hisbuf3_7[14]), .Y(n682) );
  NAND4X1 U729 ( .A(n685), .B(n684), .C(n683), .D(n682), .Y(n686) );
  AOI21X1 U730 ( .A0(n597), .A1(n687), .B0(n686), .Y(n689) );
  AOI22X1 U731 ( .A0(n657), .A1(i_hisbuf1_4[12]), .B0(n751), .B1(i_hisbuf2_5[12]), .Y(n694) );
  AOI22X1 U732 ( .A0(n640), .A1(i_hisbuf0_4[12]), .B0(n752), .B1(i_hisbuf3_3[12]), .Y(n693) );
  AOI22X1 U733 ( .A0(n753), .A1(i_hisbuf3_5[12]), .B0(n641), .B1(i_hisbuf0_6[12]), .Y(n692) );
  AOI22X1 U734 ( .A0(n642), .A1(i_hisbuf1_6[12]), .B0(n754), .B1(i_hisbuf3_6[12]), .Y(n691) );
  NAND4X1 U735 ( .A(n694), .B(n693), .C(n692), .D(n691), .Y(n700) );
  AOI22X1 U736 ( .A0(n663), .A1(i_hisbuf0_5[12]), .B0(n759), .B1(i_hisbuf3_4[12]), .Y(n698) );
  AOI22X1 U737 ( .A0(n564), .A1(i_hisbuf0_7[12]), .B0(n664), .B1(i_hisbuf1_5[12]), .Y(n697) );
  AOI22X1 U738 ( .A0(n666), .A1(i_hisbuf2_6[12]), .B0(n760), .B1(i_hisbuf2_7[12]), .Y(n696) );
  AOI22X1 U739 ( .A0(n667), .A1(i_hisbuf1_7[12]), .B0(n761), .B1(i_hisbuf3_7[12]), .Y(n695) );
  NAND4X1 U740 ( .A(n698), .B(n697), .C(n696), .D(n695), .Y(n699) );
  AOI21X1 U741 ( .A0(n597), .A1(n700), .B0(n699), .Y(n702) );
  AOI22X1 U742 ( .A0(n769), .A1(i_hisbuf2_3[12]), .B0(n732), .B1(i_agg_su_count_a[12]), .Y(n701) );
  AOI22X1 U743 ( .A0(n657), .A1(i_hisbuf1_4[9]), .B0(n751), .B1(i_hisbuf2_5[9]), .Y(n709) );
  AOI22X1 U744 ( .A0(n640), .A1(i_hisbuf0_4[9]), .B0(n704), .B1(i_hisbuf3_3[9]), .Y(n708) );
  AOI22X1 U745 ( .A0(n753), .A1(i_hisbuf3_5[9]), .B0(n641), .B1(i_hisbuf0_6[9]), .Y(n707) );
  AOI22X1 U746 ( .A0(n642), .A1(i_hisbuf1_6[9]), .B0(n705), .B1(i_hisbuf3_6[9]), .Y(n706) );
  NAND4X1 U747 ( .A(n709), .B(n708), .C(n707), .D(n706), .Y(n717) );
  AOI22X1 U748 ( .A0(n663), .A1(i_hisbuf0_5[9]), .B0(n710), .B1(i_hisbuf3_4[9]), .Y(n715) );
  AOI22X1 U749 ( .A0(n564), .A1(i_hisbuf0_7[9]), .B0(n664), .B1(i_hisbuf1_5[9]), .Y(n714) );
  AOI22X1 U750 ( .A0(n666), .A1(i_hisbuf2_6[9]), .B0(n760), .B1(i_hisbuf2_7[9]), .Y(n713) );
  AOI22X1 U751 ( .A0(n667), .A1(i_hisbuf1_7[9]), .B0(n711), .B1(i_hisbuf3_7[9]), .Y(n712) );
  NAND4X1 U752 ( .A(n715), .B(n714), .C(n713), .D(n712), .Y(n716) );
  AOI21X1 U753 ( .A0(n597), .A1(n717), .B0(n716), .Y(n719) );
  AOI22X1 U754 ( .A0(n657), .A1(i_hisbuf1_4[11]), .B0(n751), .B1(i_hisbuf2_5[11]), .Y(n724) );
  AOI22X1 U755 ( .A0(n640), .A1(i_hisbuf0_4[11]), .B0(n752), .B1(i_hisbuf3_3[11]), .Y(n723) );
  AOI22X1 U756 ( .A0(n753), .A1(i_hisbuf3_5[11]), .B0(n641), .B1(i_hisbuf0_6[11]), .Y(n722) );
  AOI22X1 U757 ( .A0(n642), .A1(i_hisbuf1_6[11]), .B0(n754), .B1(i_hisbuf3_6[11]), .Y(n721) );
  NAND4X1 U758 ( .A(n724), .B(n723), .C(n722), .D(n721), .Y(n730) );
  AOI22X1 U759 ( .A0(n663), .A1(i_hisbuf0_5[11]), .B0(n759), .B1(i_hisbuf3_4[11]), .Y(n728) );
  AOI22X1 U760 ( .A0(n564), .A1(i_hisbuf0_7[11]), .B0(n664), .B1(i_hisbuf1_5[11]), .Y(n727) );
  AOI22X1 U761 ( .A0(n666), .A1(i_hisbuf2_6[11]), .B0(n760), .B1(i_hisbuf2_7[11]), .Y(n726) );
  NAND4X1 U762 ( .A(n728), .B(n727), .C(n726), .D(n725), .Y(n729) );
  AOI21X1 U763 ( .A0(n597), .A1(n730), .B0(n729), .Y(n734) );
  AOI22X1 U764 ( .A0(n769), .A1(i_hisbuf2_3[11]), .B0(n732), .B1(i_agg_su_count_a[11]), .Y(n733) );
  AOI22X1 U765 ( .A0(n657), .A1(i_hisbuf1_4[13]), .B0(n736), .B1(i_hisbuf2_5[13]), .Y(n740) );
  AOI22X1 U766 ( .A0(n640), .A1(i_hisbuf0_4[13]), .B0(n752), .B1(i_hisbuf3_3[13]), .Y(n739) );
  AOI22X1 U767 ( .A0(n753), .A1(i_hisbuf3_5[13]), .B0(n641), .B1(i_hisbuf0_6[13]), .Y(n738) );
  AOI22X1 U768 ( .A0(n642), .A1(i_hisbuf1_6[13]), .B0(n754), .B1(i_hisbuf3_6[13]), .Y(n737) );
  NAND4X1 U769 ( .A(n740), .B(n739), .C(n738), .D(n737), .Y(n746) );
  AOI22X1 U770 ( .A0(n663), .A1(i_hisbuf0_5[13]), .B0(n759), .B1(i_hisbuf3_4[13]), .Y(n744) );
  AOI22X1 U771 ( .A0(n564), .A1(i_hisbuf0_7[13]), .B0(n664), .B1(i_hisbuf1_5[13]), .Y(n743) );
  AOI22X1 U772 ( .A0(n667), .A1(i_hisbuf1_7[13]), .B0(n761), .B1(i_hisbuf3_7[13]), .Y(n741) );
  NAND4X1 U773 ( .A(n744), .B(n743), .C(n742), .D(n741), .Y(n745) );
  AOI21X1 U774 ( .A0(n597), .A1(n746), .B0(n745), .Y(n748) );
  AOI22X1 U775 ( .A0(n769), .A1(i_hisbuf2_3[13]), .B0(n768), .B1(i_agg_su_count_a[13]), .Y(n747) );
  AOI22X1 U776 ( .A0(n640), .A1(i_hisbuf0_4[10]), .B0(n752), .B1(i_hisbuf3_3[10]), .Y(n757) );
  AOI22X1 U777 ( .A0(n753), .A1(i_hisbuf3_5[10]), .B0(n641), .B1(i_hisbuf0_6[10]), .Y(n756) );
  AOI22X1 U778 ( .A0(n642), .A1(i_hisbuf1_6[10]), .B0(n754), .B1(i_hisbuf3_6[10]), .Y(n755) );
  NAND4X1 U779 ( .A(n758), .B(n757), .C(n756), .D(n755), .Y(n767) );
  AOI22X1 U780 ( .A0(n663), .A1(i_hisbuf0_5[10]), .B0(n759), .B1(i_hisbuf3_4[10]), .Y(n765) );
  AOI22X1 U781 ( .A0(n564), .A1(i_hisbuf0_7[10]), .B0(n664), .B1(i_hisbuf1_5[10]), .Y(n764) );
  AOI22X1 U782 ( .A0(n666), .A1(i_hisbuf2_6[10]), .B0(n760), .B1(i_hisbuf2_7[10]), .Y(n763) );
  AOI22X1 U783 ( .A0(n667), .A1(i_hisbuf1_7[10]), .B0(n761), .B1(i_hisbuf3_7[10]), .Y(n762) );
  NAND4X1 U784 ( .A(n765), .B(n764), .C(n763), .D(n762), .Y(n766) );
  AOI21X1 U785 ( .A0(n597), .A1(n767), .B0(n766), .Y(n771) );
  AOI22X1 U786 ( .A0(n769), .A1(i_hisbuf2_3[10]), .B0(n768), .B1(i_agg_su_count_a[10]), .Y(n770) );
  AOI22X1 U787 ( .A0(n170), .A1(i_hisbuf0_3[23]), .B0(n168), .B1(i_hisbuf0_2[23]), .Y(n782) );
  AOI22X1 U788 ( .A0(n814), .A1(i_hisbuf2_2[23]), .B0(i_hisbuf1_2[23]), .B1(n166), .Y(n781) );
  AOI22X1 U789 ( .A0(n838), .A1(i_hisbuf1_0[23]), .B0(i_hisbuf2_0[23]), .B1(n830), .Y(n776) );
  AOI22X1 U790 ( .A0(n815), .A1(i_hisbuf3_0[23]), .B0(n836), .B1(i_hisbuf2_1[23]), .Y(n775) );
  AOI22X1 U791 ( .A0(n843), .A1(i_hisbuf3_1[23]), .B0(n130), .B1(i_spare_config[23]), .Y(n773) );
  NAND4X1 U792 ( .A(n776), .B(n775), .C(n774), .D(n773), .Y(n779) );
  AOI22X1 U793 ( .A0(n165), .A1(i_hisbuf1_3[23]), .B0(n807), .B1(i_hisbuf3_2[23]), .Y(n777) );
  AO21X1 U794 ( .A0(n823), .A1(i_hisbuf0_0[23]), .B0(n777_inv), .Y(n778) );
  AOI22X1 U795 ( .A0(n170), .A1(i_hisbuf0_3[18]), .B0(n168), .B1(i_hisbuf0_2[18]), .Y(n792) );
  AOI22X1 U796 ( .A0(n814), .A1(i_hisbuf2_2[18]), .B0(i_hisbuf1_2[18]), .B1(n166), .Y(n791) );
  AOI22X1 U797 ( .A0(n838), .A1(i_hisbuf1_0[18]), .B0(i_hisbuf2_0[18]), .B1(n830), .Y(n786) );
  AOI22X1 U798 ( .A0(n815), .A1(i_hisbuf3_0[18]), .B0(n836), .B1(i_hisbuf2_1[18]), .Y(n785) );
  AOI22X1 U799 ( .A0(n311), .A1(i_hisbuf0_1[18]), .B0(n816), .B1(i_hisbuf1_1[18]), .Y(n784) );
  AOI22X1 U800 ( .A0(n843), .A1(i_hisbuf3_1[18]), .B0(n130), .B1(i_spare_config[18]), .Y(n783) );
  NAND4X1 U801 ( .A(n786), .B(n785), .C(n784), .D(n783), .Y(n789) );
  AOI22X1 U802 ( .A0(n165), .A1(i_hisbuf1_3[18]), .B0(n821), .B1(i_hisbuf3_2[18]), .Y(n787) );
  AO21X1 U803 ( .A0(n823), .A1(i_hisbuf0_0[18]), .B0(n787_inv), .Y(n788) );
  AOI22X1 U804 ( .A0(n170), .A1(i_hisbuf0_3[19]), .B0(n168), .B1(i_hisbuf0_2[19]), .Y(n802) );
  AOI22X1 U805 ( .A0(n814), .A1(i_hisbuf2_2[19]), .B0(i_hisbuf1_2[19]), .B1(n166), .Y(n801) );
  AOI22X1 U806 ( .A0(n838), .A1(i_hisbuf1_0[19]), .B0(i_hisbuf2_0[19]), .B1(n830), .Y(n796) );
  AOI22X1 U807 ( .A0(n815), .A1(i_hisbuf3_0[19]), .B0(n836), .B1(i_hisbuf2_1[19]), .Y(n795) );
  AOI22X1 U808 ( .A0(n311), .A1(i_hisbuf0_1[19]), .B0(n816), .B1(i_hisbuf1_1[19]), .Y(n794) );
  AOI22X1 U809 ( .A0(n843), .A1(i_hisbuf3_1[19]), .B0(n130), .B1(i_spare_config[19]), .Y(n793) );
  NAND4X1 U810 ( .A(n796), .B(n795), .C(n794), .D(n793), .Y(n799) );
  AOI22X1 U811 ( .A0(n165), .A1(i_hisbuf1_3[19]), .B0(n807), .B1(i_hisbuf3_2[19]), .Y(n797) );
  AO21X1 U812 ( .A0(n823), .A1(i_hisbuf0_0[19]), .B0(n797_inv), .Y(n798) );
  AOI21X1 U813 ( .A0(n852), .A1(n799), .B0(n798), .Y(n800) );
  AOI22X1 U814 ( .A0(n170), .A1(i_hisbuf0_3[20]), .B0(n168), .B1(i_hisbuf0_2[20]), .Y(n813) );
  AOI22X1 U815 ( .A0(n814), .A1(i_hisbuf2_2[20]), .B0(i_hisbuf1_2[20]), .B1(n166), .Y(n812) );
  AOI22X1 U816 ( .A0(n838), .A1(i_hisbuf1_0[20]), .B0(i_hisbuf2_0[20]), .B1(n830), .Y(n806) );
  AOI22X1 U817 ( .A0(n311), .A1(i_hisbuf0_1[20]), .B0(n816), .B1(i_hisbuf1_1[20]), .Y(n804) );
  AOI22X1 U818 ( .A0(n843), .A1(i_hisbuf3_1[20]), .B0(n130), .B1(i_spare_config[20]), .Y(n803) );
  NAND4X1 U819 ( .A(n806), .B(n805), .C(n804), .D(n803), .Y(n810) );
  AOI22X1 U820 ( .A0(n165), .A1(i_hisbuf1_3[20]), .B0(n807), .B1(i_hisbuf3_2[20]), .Y(n808) );
  AO21X1 U821 ( .A0(n823), .A1(i_hisbuf0_0[20]), .B0(n808_inv), .Y(n809) );
  AOI21X1 U822 ( .A0(n852), .A1(n810), .B0(n809), .Y(n811) );
  AOI22X1 U823 ( .A0(n170), .A1(i_hisbuf0_3[16]), .B0(n168), .B1(i_hisbuf0_2[16]), .Y(n828) );
  AOI22X1 U824 ( .A0(n814), .A1(i_hisbuf2_2[16]), .B0(i_hisbuf1_2[16]), .B1(n166), .Y(n827) );
  AOI22X1 U825 ( .A0(n838), .A1(i_hisbuf1_0[16]), .B0(i_hisbuf2_0[16]), .B1(n830), .Y(n820) );
  AOI22X1 U826 ( .A0(n815), .A1(i_hisbuf3_0[16]), .B0(n836), .B1(i_hisbuf2_1[16]), .Y(n819) );
  AOI22X1 U827 ( .A0(n311), .A1(i_hisbuf0_1[16]), .B0(n816), .B1(i_hisbuf1_1[16]), .Y(n818) );
  AOI22X1 U828 ( .A0(n843), .A1(i_hisbuf3_1[16]), .B0(n130), .B1(i_spare_config[16]), .Y(n817) );
  NAND4X1 U829 ( .A(n820), .B(n819), .C(n818), .D(n817), .Y(n825) );
  AOI22X1 U830 ( .A0(n165), .A1(i_hisbuf1_3[16]), .B0(n821), .B1(i_hisbuf3_2[16]), .Y(n822) );
  AO21X1 U831 ( .A0(n823), .A1(i_hisbuf0_0[16]), .B0(n822_inv), .Y(n824) );
  AOI21X1 U832 ( .A0(n852), .A1(n825), .B0(n824), .Y(n826) );
  INVX2 U833 ( .A(scan_iso_or7), .Y(n835) );
  AOI22X1 U834 ( .A0(n830), .A1(i_hisbuf2_0[0]), .B0(n829), .B1(o_dbg_config[0]), .Y(n833) );
  AOI22X1 U835 ( .A0(n831), .A1(i_hisbuf1_2[0]), .B0(n130), .B1(i_spare_config[0]), .Y(n832) );
  OAI211X1 U836 ( .A0(n835), .A1(n834), .B0(n833), .C0(n832), .Y(n855) );
  AOI22X1 U837 ( .A0(n837), .A1(i_hisbuf3_0[0]), .B0(n836), .B1(i_hisbuf2_1[0]), .Y(n841) );
  NAND2X1 U838 ( .A(n841), .B(n840), .Y(n854) );
  AOI22X1 U839 ( .A0(n816), .A1(i_hisbuf1_1[0]), .B0(n843), .B1(i_hisbuf3_1[0]), .Y(n851) );
  AOI22X1 U840 ( .A0(n159), .A1(i_hisbuf0_0[0]), .B0(n311), .B1(i_hisbuf0_1[0]), .Y(n850) );
  AOI22X1 U841 ( .A0(n845), .A1(i_hisbuf3_2[0]), .B0(n844), .B1(i_hisbuf0_2[0]), .Y(n849) );
  AOI22X1 U842 ( .A0(n847), .A1(i_hisbuf0_3[0]), .B0(n846), .B1(i_hisbuf1_3[0]), .Y(n848) );
  NAND4X1 U843 ( .A(n851), .B(n850), .C(n849), .D(n848), .Y(n853));
  OAI31X1 U844 ( .A0(n855), .A1(n854), .A2(n853), .B0(n852), .Y(n856) );
  AO21X1 U845 ( .A0(n857), .A1(i_hisbuf2_2[0]), .B0(n856_inv), .Y(N422) );
  INVX1 U186_INV ( .A(n353), .Y(n353_inv) );
  INVX1 U264_INV ( .A(n188), .Y(n188_inv) );
  INVX1 U274_INV ( .A(n199), .Y(n199_inv) );
  INVX1 U434_INV ( .A(n343), .Y(n343_inv) );
  INVX1 U453_INV ( .A(n363), .Y(n363_inv) );
  INVX1 U794_INV ( .A(n777), .Y(n777_inv) );
  INVX1 U803_INV ( .A(n787), .Y(n787_inv) );
  INVX1 U812_INV ( .A(n797), .Y(n797_inv) );
  INVX1 U821_INV ( .A(n808), .Y(n808_inv) );
  INVX1 U831_INV ( .A(n822), .Y(n822_inv) );
  INVX1 U845_INV ( .A(n856), .Y(n856_inv) );
  survik u_survik ( .clk(clk), .i_reset_(n128), 
 .i_sw_init(1'b0), .o_spare_config(o_spare_config), .o_adj_config(
 o_adj_config), .o_dbg_config(o_dbg_config[0]), .w_load_spare_config(
 w_load_spare_config), .w_load_adj_config(w_load_adj_config), 
 .w_load_dbg_config(w_load_dbg_config), .f32_data({n_94_, n_95_, n_96_, 
 n_97_, n_98_, n_99_, n_100_, n_101_, n_102_, n_103_, n_104_, n_105_, 
 n_106_, n_107_, n_108_, n_109_, n_110_, n_111_, n_112_, n_113_, n_114_, 
 test_so1, n_116_, n_117_, n_118_, n_119_, n_120_, n_121_, n_122_, 
 n_123_, n_124_, n_125_}), .scan_iso_or(scan_iso_or6), .test_se(test_se), .scan_iso_or1(scan_iso_or7), .scan_iso_or2(scan_iso_or8), .scan_iso_or3(
 scan_iso_or9), .test_si(o_reg_read), .scan_enable(scan_enable) );
  TLATNTSCAX12 clk_gate_mux ( .CK(clk), .E(N421), .ECK(net121966),  .SE(scan_enable) );
  TLATNTSCAX12 clk_gate_addr ( .CK(clk), .E(N410), .ECK(net121972),  .SE(scan_enable) );
  TLATNTSCAX12 clk_gate_data ( .CK(clk), .E(i_wr_strb), .ECK(net121977),  .SE( scan_enable) );
  NAND2BX1 U43 ( .AN(scan_iso_or3), .B(scan_iso_or4), .Y(n386) );
  INVX4 U12 ( .A(n131), .Y(n500) );
  OR2X1 U27 ( .A(n379), .B(n500), .Y(n381) );
  NOR2BX2 U202 ( .AN(n836), .B(n132), .Y(n134) );
  NOR2BX2 U204 ( .AN(n843), .B(n132), .Y(n328) );
  NOR2X4 U25 ( .A(n834), .B(n395), .Y(n564) );
  INVX2 U14 ( .A(n126), .Y(n127) );
  INVX4 U13 ( .A(i_reset_), .Y(n126) );
  NOR3X2 U3 ( .A(n379), .B(n393), .C(n500), .Y(n750) );
  INVX4 U4 ( .A(n852), .Y(n132) );
  NOR2X2 U20 ( .A(n158), .B(f_ack), .Y(n335) );
  BUFX2 U21 ( .A(n837), .Y(n815) );
  NAND3X1 U32 ( .A(n370), .B(n372), .C(scan_iso_or1), .Y(n379) );
  NAND3X2 U53 ( .A(n371), .B(n370), .C(scan_iso_or), .Y(n169) );
  INVX8 U74 ( .A(n126), .Y(n128) );
  AND2X1 o_reg_addr_reg_6__scan_iso_or ( .A(o_reg_addr[6]), .B(test_se), .Y(scan_iso_or) );
  AND2X1 o_reg_addr_reg_5__scan_iso_or ( .A(o_reg_addr[5]), .B(test_se), .Y(scan_iso_or1) );
  AND2X1 o_reg_addr_reg_4__scan_iso_or ( .A(o_reg_addr[4]), .B(test_se), .Y(scan_iso_or2) );
  AND2X1 o_reg_addr_reg_3__scan_iso_or ( .A(o_reg_addr[3]), .B(test_se), .Y(scan_iso_or3) );
  AND2X1 o_reg_addr_reg_2__scan_iso_or ( .A(o_reg_addr[2]), .B(test_se), .Y(scan_iso_or4) );
  AND2X1 o_reg_addr_reg_7__scan_iso_or ( .A(o_reg_addr[7]), .B(test_se), .Y(scan_iso_or5) );
  AND2X1 o_reg_addr_reg_1__scan_iso_or ( .A(n862), .B(test_se), .Y(o_reg_addr_reg_1__scan_iso_or_n) );
  AND2X1 o_reg_addr_reg_0__scan_iso_or ( .A(n863), .B(test_se), .Y(o_reg_addr_reg_0__scan_iso_or_n) );
  MX2X2 f32_data_reg_11__ti_over_mux ( .A(n_113_), .B(test_si1), .S0(raw_scan_en), .Y(n1) );
endmodule
module survik (clk, i_reset_, i_sw_init, o_spare_config, 
 o_adj_config, o_dbg_config, w_load_spare_config, w_load_adj_config, 
 w_load_dbg_config, f32_data, scan_iso_or, test_se, scan_iso_or1, 
 scan_iso_or2, scan_iso_or3, test_si, scan_enable);
  output [31:0] o_spare_config;
  output [15:0] o_adj_config;
  output [0:0] o_dbg_config;
  input [31:0] f32_data;
  input clk, i_reset_, i_sw_init, w_load_spare_config, w_load_adj_config,
 w_load_dbg_config, test_se, test_si, scan_enable;
  output scan_iso_or, scan_iso_or1, scan_iso_or2, scan_iso_or3;
  wire net121994, net122000, n37, n38, n39, n51;

  SDFFRX1 o_dbg_config_reg_0_ ( .D(n51), .SI(o_adj_config[15]), .SE(scan_enable), .CK(clk), .RN(n39), .Q(o_dbg_config[0]) );
  SDFFRX1 o_spare_config_reg_31_ ( .D(f32_data[31]), .SI(o_spare_config[30]), .SE(scan_enable), .CK(net121994), .RN(n38),  .Q(o_spare_config[31]) );
  SDFFRX1 o_spare_config_reg_30_ ( .D(f32_data[30]), .SI(o_spare_config[29]), .SE(scan_enable), .CK(net121994), .RN(n38),  .Q(o_spare_config[30]) );
  SDFFRX1 o_spare_config_reg_29_ ( .D(f32_data[29]), .SI(o_spare_config[28]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[29]) );
  SDFFRX1 o_spare_config_reg_28_ ( .D(f32_data[28]), .SI(o_spare_config[27]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[28]) );
  SDFFRX1 o_spare_config_reg_27_ ( .D(f32_data[27]), .SI(o_spare_config[26]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[27]) );
  SDFFRX1 o_spare_config_reg_26_ ( .D(f32_data[26]), .SI(o_spare_config[25]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[26]) );
  SDFFRX1 o_spare_config_reg_25_ ( .D(f32_data[25]), .SI(o_spare_config[24]), .SE(scan_enable), .CK(net121994), .RN(n38),  .Q(o_spare_config[25]) );
  SDFFRX1 o_spare_config_reg_24_ ( .D(f32_data[24]), .SI(o_spare_config[23]), .SE(scan_enable), .CK(net121994), .RN(n38),  .Q(o_spare_config[24]) );
  SDFFRX1 o_spare_config_reg_23_ ( .D(f32_data[23]), .SI(o_spare_config[22]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[23]) );
  SDFFRX1 o_spare_config_reg_22_ ( .D(f32_data[22]), .SI(o_spare_config[21]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[22]) );
  SDFFRX1 o_spare_config_reg_21_ ( .D(f32_data[21]), .SI(o_spare_config[20]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[21]) );
  SDFFRX1 o_spare_config_reg_20_ ( .D(f32_data[20]), .SI(o_spare_config[19]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[20]) );
  SDFFRX1 o_spare_config_reg_19_ ( .D(f32_data[19]), .SI(o_spare_config[18]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[19]) );
  SDFFRX1 o_spare_config_reg_18_ ( .D(f32_data[18]), .SI(o_spare_config[17]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[18]) );
  SDFFRX1 o_spare_config_reg_17_ ( .D(f32_data[17]), .SI(o_spare_config[16]), .SE(scan_enable), .CK(net121994), .RN(n38),  .Q(o_spare_config[17]) );
  SDFFRX1 o_spare_config_reg_16_ ( .D(f32_data[16]), .SI(o_spare_config[15]), .SE(scan_enable), .CK(net121994), .RN(n38),  .Q(o_spare_config[16]) );
  SDFFRX1 o_spare_config_reg_15_ ( .D(f32_data[15]), .SI(o_spare_config[14]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[15]) );
  SDFFRX1 o_spare_config_reg_14_ ( .D(f32_data[14]), .SI(o_spare_config[13]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[14]) );
  SDFFRX1 o_spare_config_reg_13_ ( .D(f32_data[13]), .SI(o_spare_config[12]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[13]) );
  SDFFRX1 o_spare_config_reg_12_ ( .D(f32_data[12]), .SI(o_spare_config[11]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[12]) );
  SDFFRX1 o_spare_config_reg_11_ ( .D(f32_data[11]), .SI(o_spare_config[10]), .SE(scan_enable), .CK(net121994), .RN(n38),  .Q(o_spare_config[11]) );
  SDFFRX1 o_spare_config_reg_10_ ( .D(f32_data[10]), .SI(o_spare_config[9]), .SE(scan_enable), .CK(net121994), .RN(n38),  .Q(o_spare_config[10]) );
  SDFFRX1 o_spare_config_reg_9_ ( .D(f32_data[9]), .SI(o_spare_config[8]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[9]) );
  SDFFRX1 o_spare_config_reg_8_ ( .D(f32_data[8]), .SI(o_spare_config[7]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[8]) );
  SDFFRX1 o_spare_config_reg_7_ ( .D(f32_data[7]), .SI(o_spare_config[6]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[7]) );
  SDFFRX1 o_spare_config_reg_6_ ( .D(f32_data[6]), .SI(o_spare_config[5]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[6]) );
  SDFFRX1 o_spare_config_reg_5_ ( .D(f32_data[5]), .SI(o_spare_config[4]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[5]) );
  SDFFRX1 o_spare_config_reg_4_ ( .D(f32_data[4]), .SI(o_spare_config[3]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[4]) );
  SDFFRX1 o_spare_config_reg_3_ ( .D(f32_data[3]), .SI(o_spare_config[2]), .SE(scan_enable), .CK(net121994), .RN(n39),  .Q(o_spare_config[3]) );
  SDFFRX1 o_spare_config_reg_2_ ( .D(f32_data[2]), .SI(o_spare_config[1]), .SE(scan_enable), .CK(net121994), .RN(n38),  .Q(o_spare_config[2]) );
  SDFFRX1 o_spare_config_reg_1_ ( .D(f32_data[1]), .SI(o_spare_config[0]), .SE(scan_enable), .CK(net121994), .RN(n38),  .Q(o_spare_config[1]) );
  SDFFRX1 o_spare_config_reg_0_ ( .D(f32_data[0]), .SI(o_dbg_config[0]), .SE(scan_enable), .CK(net121994), .RN(n38), .Q(o_spare_config[0]) );
  SDFFRX1 o_adj_config_reg_15_ ( .D(f32_data[15]), .SI(o_adj_config[14]), .SE(scan_enable), .CK(net122000), .RN(n38),  .Q(o_adj_config[15]) );
  SDFFRX1 o_adj_config_reg_14_ ( .D(f32_data[14]), .SI(o_adj_config[13]), .SE(scan_enable), .CK(net122000), .RN(n38),  .Q(o_adj_config[14]) );
  SDFFRX1 o_adj_config_reg_13_ ( .D(f32_data[13]), .SI(o_adj_config[12]), .SE(scan_enable), .CK(net122000), .RN(n38),  .Q(o_adj_config[13]) );
  SDFFRX1 o_adj_config_reg_12_ ( .D(f32_data[12]), .SI(o_adj_config[11]), .SE(scan_enable), .CK(net122000), .RN(n38),  .Q(o_adj_config[12]) );
  SDFFRX1 o_adj_config_reg_11_ ( .D(f32_data[11]), .SI(o_adj_config[10]), .SE(scan_enable), .CK(net122000), .RN(n39),  .Q(o_adj_config[11]) );
  SDFFRX1 o_adj_config_reg_10_ ( .D(f32_data[10]), .SI(o_adj_config[9]), .SE(scan_enable), .CK(net122000), .RN(i_reset_), .Q(o_adj_config[10]) );
  SDFFRX1 o_adj_config_reg_9_ ( .D(f32_data[9]), .SI(o_adj_config[8]), .SE(scan_enable), .CK(net122000), .RN(i_reset_), .Q(o_adj_config[9]) );
  SDFFRX1 o_adj_config_reg_8_ ( .D(f32_data[8]), .SI(o_adj_config[7]), .SE(scan_enable), .CK(net122000), .RN(i_reset_), .Q(o_adj_config[8]) );
  SDFFRX1 o_adj_config_reg_7_ ( .D(f32_data[7]), .SI(o_adj_config[6]), .SE(scan_enable), .CK(net122000), .RN(i_reset_), .Q(o_adj_config[7]) );
  SDFFRX1 o_adj_config_reg_6_ ( .D(f32_data[6]), .SI(o_adj_config[5]), .SE(scan_enable), .CK(net122000), .RN(i_reset_), .Q(o_adj_config[6]) );
  SDFFRX1 o_adj_config_reg_5_ ( .D(f32_data[5]), .SI(o_adj_config[4]), .SE(scan_enable), .CK(net122000), .RN(i_reset_), .Q(o_adj_config[5]) );
  SDFFRX1 o_adj_config_reg_4_ ( .D(f32_data[4]), .SI(o_adj_config[3]), .SE(scan_enable), .CK(net122000), .RN(i_reset_), .Q(o_adj_config[4]) );
  SDFFRX1 o_adj_config_reg_3_ ( .D(f32_data[3]), .SI(o_adj_config[2]), .SE(scan_enable), .CK(net122000), .RN(i_reset_), .Q(o_adj_config[3]) );
  SDFFRX1 o_adj_config_reg_2_ ( .D(f32_data[2]), .SI(o_adj_config[1]), .SE(scan_enable), .CK(net122000), .RN(i_reset_), .Q(o_adj_config[2]) );
  SDFFRX1 o_adj_config_reg_1_ ( .D(f32_data[1]), .SI(o_adj_config[0]), .SE(scan_enable), .CK(net122000), .RN(i_reset_), .Q(o_adj_config[1]) );
  SDFFRX1 o_adj_config_reg_0_ ( .D(f32_data[0]), .SI(test_si), .SE(scan_enable), .CK(net122000), .RN(i_reset_), .Q(o_adj_config[0]) );
  MX2X1 U7 ( .A(o_dbg_config[0]), .B(f32_data[0]), .S0(w_load_dbg_config), .Y(n51) );
  TLATNTSCAX12 clk_gate_spare_config ( .CK(clk), .E(w_load_spare_config), .ECK(net121994), .SE(scan_enable) );
  TLATNTSCAX12 clk_gate_config ( .CK(clk), .E(w_load_adj_config), .ECK(net122000), .SE(scan_enable) );
  INVX2 U4 ( .A(i_reset_), .Y(n37) );
  BUFX8 U3 ( .A(i_reset_), .Y(n39) );
  INVX6 U5 ( .A(n37), .Y(n38) );
  AND2X1 o_adj_config_reg_1__scan_iso_or ( .A(o_adj_config[1]), .B(test_se), .Y(scan_iso_or) );
  AND2X1 o_adj_config_reg_0__scan_iso_or ( .A(o_adj_config[0]), .B(test_se), .Y(scan_iso_or1) );
  AND2X1 o_adj_config_reg_2__scan_iso_or ( .A(o_adj_config[2]), .B(test_se), .Y(scan_iso_or2) );
  AND2X1 o_adj_config_reg_3__scan_iso_or ( .A(o_adj_config[3]), .B(test_se), .Y(scan_iso_or3) );
endmodule
